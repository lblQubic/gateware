assign dspif.weight_bias[0][0]= dspregs.W_Q0_0_0_0;
assign dspif.weight_bias[0][1]= dspregs.W_Q0_0_0_1;
assign dspif.weight_bias[0][2]= dspregs.W_Q0_0_0_2;
assign dspif.weight_bias[0][3]= dspregs.W_Q0_0_0_3;
assign dspif.weight_bias[0][4]= dspregs.W_Q0_0_0_4;
assign dspif.weight_bias[0][5]= dspregs.W_Q0_0_0_5;
assign dspif.weight_bias[0][6]= dspregs.W_Q0_0_0_6;
assign dspif.weight_bias[0][7]= dspregs.W_Q0_0_0_7;
assign dspif.weight_bias[0][8]= dspregs.W_Q0_0_1_0;
assign dspif.weight_bias[0][9]= dspregs.W_Q0_0_1_1;
assign dspif.weight_bias[0][10]=dspregs.W_Q0_0_1_2;
assign dspif.weight_bias[0][11]=dspregs.W_Q0_0_1_3;
assign dspif.weight_bias[0][12]=dspregs.W_Q0_0_1_4;
assign dspif.weight_bias[0][13]=dspregs.W_Q0_0_1_5;
assign dspif.weight_bias[0][14]=dspregs.W_Q0_0_1_6;
assign dspif.weight_bias[0][15]=dspregs.W_Q0_0_1_7;
assign dspif.weight_bias[0][16]=dspregs.W_Q0_1_0_0;
assign dspif.weight_bias[0][17]=dspregs.W_Q0_1_0_1;
assign dspif.weight_bias[0][18]=dspregs.W_Q0_1_0_2;
assign dspif.weight_bias[0][19]=dspregs.W_Q0_1_0_3;
assign dspif.weight_bias[0][20]=dspregs.W_Q0_1_1_0;
assign dspif.weight_bias[0][21]=dspregs.W_Q0_1_1_1;
assign dspif.weight_bias[0][22]=dspregs.W_Q0_1_1_2;
assign dspif.weight_bias[0][23]=dspregs.W_Q0_1_1_3;
assign dspif.weight_bias[0][24]=dspregs.W_Q0_1_2_0;
assign dspif.weight_bias[0][25]=dspregs.W_Q0_1_2_1;
assign dspif.weight_bias[0][26]=dspregs.W_Q0_1_2_2;
assign dspif.weight_bias[0][27]=dspregs.W_Q0_1_2_3;
assign dspif.weight_bias[0][28]=dspregs.W_Q0_1_3_0;
assign dspif.weight_bias[0][29]=dspregs.W_Q0_1_3_1;
assign dspif.weight_bias[0][30]=dspregs.W_Q0_1_3_2;
assign dspif.weight_bias[0][31]=dspregs.W_Q0_1_3_3;
assign dspif.weight_bias[0][32]=dspregs.W_Q0_1_4_0;
assign dspif.weight_bias[0][33]=dspregs.W_Q0_1_4_1;
assign dspif.weight_bias[0][34]=dspregs.W_Q0_1_4_2;
assign dspif.weight_bias[0][35]=dspregs.W_Q0_1_4_3;
assign dspif.weight_bias[0][36]=dspregs.W_Q0_1_5_0;
assign dspif.weight_bias[0][37]=dspregs.W_Q0_1_5_1;
assign dspif.weight_bias[0][38]=dspregs.W_Q0_1_5_2;
assign dspif.weight_bias[0][39]=dspregs.W_Q0_1_5_3;
assign dspif.weight_bias[0][40]=dspregs.W_Q0_1_6_0;
assign dspif.weight_bias[0][41]=dspregs.W_Q0_1_6_1;
assign dspif.weight_bias[0][42]=dspregs.W_Q0_1_6_2;
assign dspif.weight_bias[0][43]=dspregs.W_Q0_1_6_3;
assign dspif.weight_bias[0][44]=dspregs.W_Q0_1_7_0;
assign dspif.weight_bias[0][45]=dspregs.W_Q0_1_7_1;
assign dspif.weight_bias[0][46]=dspregs.W_Q0_1_7_2;
assign dspif.weight_bias[0][47]=dspregs.W_Q0_1_7_3;
assign dspif.weight_bias[0][48]=dspregs.W_Q0_2_0_0;
assign dspif.weight_bias[0][49]=dspregs.W_Q0_2_1_0;
assign dspif.weight_bias[0][50]=dspregs.W_Q0_2_2_0;
assign dspif.weight_bias[0][51]=dspregs.W_Q0_2_3_0;
assign dspif.weight_bias[0][52]=dspregs.B_Q0_0_0;
assign dspif.weight_bias[0][53]=dspregs.B_Q0_0_1;
assign dspif.weight_bias[0][54]=dspregs.B_Q0_0_2;
assign dspif.weight_bias[0][55]=dspregs.B_Q0_0_3;
assign dspif.weight_bias[0][56]=dspregs.B_Q0_0_4;
assign dspif.weight_bias[0][57]=dspregs.B_Q0_0_5;
assign dspif.weight_bias[0][58]=dspregs.B_Q0_0_6;
assign dspif.weight_bias[0][59]=dspregs.B_Q0_0_7;
assign dspif.weight_bias[0][60]=dspregs.B_Q0_1_0;
assign dspif.weight_bias[0][61]=dspregs.B_Q0_1_1;
assign dspif.weight_bias[0][62]=dspregs.B_Q0_1_2;
assign dspif.weight_bias[0][63]=dspregs.B_Q0_1_3;
assign dspif.weight_bias[0][64]=dspregs.B_Q0_2_0;
assign dspif.weight_bias[1][0]= dspregs.W_Q1_0_0_0;
assign dspif.weight_bias[1][1]= dspregs.W_Q1_0_0_1;
assign dspif.weight_bias[1][2]= dspregs.W_Q1_0_0_2;
assign dspif.weight_bias[1][3]= dspregs.W_Q1_0_0_3;
assign dspif.weight_bias[1][4]= dspregs.W_Q1_0_0_4;
assign dspif.weight_bias[1][5]= dspregs.W_Q1_0_0_5;
assign dspif.weight_bias[1][6]= dspregs.W_Q1_0_0_6;
assign dspif.weight_bias[1][7]= dspregs.W_Q1_0_0_7;
assign dspif.weight_bias[1][8]= dspregs.W_Q1_0_1_0;
assign dspif.weight_bias[1][9]= dspregs.W_Q1_0_1_1;
assign dspif.weight_bias[1][10]=dspregs.W_Q1_0_1_2;
assign dspif.weight_bias[1][11]=dspregs.W_Q1_0_1_3;
assign dspif.weight_bias[1][12]=dspregs.W_Q1_0_1_4;
assign dspif.weight_bias[1][13]=dspregs.W_Q1_0_1_5;
assign dspif.weight_bias[1][14]=dspregs.W_Q1_0_1_6;
assign dspif.weight_bias[1][15]=dspregs.W_Q1_0_1_7;
assign dspif.weight_bias[1][16]=dspregs.W_Q1_1_0_0;
assign dspif.weight_bias[1][17]=dspregs.W_Q1_1_0_1;
assign dspif.weight_bias[1][18]=dspregs.W_Q1_1_0_2;
assign dspif.weight_bias[1][19]=dspregs.W_Q1_1_0_3;
assign dspif.weight_bias[1][20]=dspregs.W_Q1_1_1_0;
assign dspif.weight_bias[1][21]=dspregs.W_Q1_1_1_1;
assign dspif.weight_bias[1][22]=dspregs.W_Q1_1_1_2;
assign dspif.weight_bias[1][23]=dspregs.W_Q1_1_1_3;
assign dspif.weight_bias[1][24]=dspregs.W_Q1_1_2_0;
assign dspif.weight_bias[1][25]=dspregs.W_Q1_1_2_1;
assign dspif.weight_bias[1][26]=dspregs.W_Q1_1_2_2;
assign dspif.weight_bias[1][27]=dspregs.W_Q1_1_2_3;
assign dspif.weight_bias[1][28]=dspregs.W_Q1_1_3_0;
assign dspif.weight_bias[1][29]=dspregs.W_Q1_1_3_1;
assign dspif.weight_bias[1][30]=dspregs.W_Q1_1_3_2;
assign dspif.weight_bias[1][31]=dspregs.W_Q1_1_3_3;
assign dspif.weight_bias[1][32]=dspregs.W_Q1_1_4_0;
assign dspif.weight_bias[1][33]=dspregs.W_Q1_1_4_1;
assign dspif.weight_bias[1][34]=dspregs.W_Q1_1_4_2;
assign dspif.weight_bias[1][35]=dspregs.W_Q1_1_4_3;
assign dspif.weight_bias[1][36]=dspregs.W_Q1_1_5_0;
assign dspif.weight_bias[1][37]=dspregs.W_Q1_1_5_1;
assign dspif.weight_bias[1][38]=dspregs.W_Q1_1_5_2;
assign dspif.weight_bias[1][39]=dspregs.W_Q1_1_5_3;
assign dspif.weight_bias[1][40]=dspregs.W_Q1_1_6_0;
assign dspif.weight_bias[1][41]=dspregs.W_Q1_1_6_1;
assign dspif.weight_bias[1][42]=dspregs.W_Q1_1_6_2;
assign dspif.weight_bias[1][43]=dspregs.W_Q1_1_6_3;
assign dspif.weight_bias[1][44]=dspregs.W_Q1_1_7_0;
assign dspif.weight_bias[1][45]=dspregs.W_Q1_1_7_1;
assign dspif.weight_bias[1][46]=dspregs.W_Q1_1_7_2;
assign dspif.weight_bias[1][47]=dspregs.W_Q1_1_7_3;
assign dspif.weight_bias[1][48]=dspregs.W_Q1_2_0_0;
assign dspif.weight_bias[1][49]=dspregs.W_Q1_2_1_0;
assign dspif.weight_bias[1][50]=dspregs.W_Q1_2_2_0;
assign dspif.weight_bias[1][51]=dspregs.W_Q1_2_3_0;
assign dspif.weight_bias[1][52]=dspregs.B_Q1_0_0;
assign dspif.weight_bias[1][53]=dspregs.B_Q1_0_1;
assign dspif.weight_bias[1][54]=dspregs.B_Q1_0_2;
assign dspif.weight_bias[1][55]=dspregs.B_Q1_0_3;
assign dspif.weight_bias[1][56]=dspregs.B_Q1_0_4;
assign dspif.weight_bias[1][57]=dspregs.B_Q1_0_5;
assign dspif.weight_bias[1][58]=dspregs.B_Q1_0_6;
assign dspif.weight_bias[1][59]=dspregs.B_Q1_0_7;
assign dspif.weight_bias[1][60]=dspregs.B_Q1_1_0;
assign dspif.weight_bias[1][61]=dspregs.B_Q1_1_1;
assign dspif.weight_bias[1][62]=dspregs.B_Q1_1_2;
assign dspif.weight_bias[1][63]=dspregs.B_Q1_1_3;
assign dspif.weight_bias[1][64]=dspregs.B_Q1_2_0;
assign dspif.weight_bias[2][0]= dspregs.W_Q2_0_0_0;
assign dspif.weight_bias[2][1]= dspregs.W_Q2_0_0_1;
assign dspif.weight_bias[2][2]= dspregs.W_Q2_0_0_2;
assign dspif.weight_bias[2][3]= dspregs.W_Q2_0_0_3;
assign dspif.weight_bias[2][4]= dspregs.W_Q2_0_0_4;
assign dspif.weight_bias[2][5]= dspregs.W_Q2_0_0_5;
assign dspif.weight_bias[2][6]= dspregs.W_Q2_0_0_6;
assign dspif.weight_bias[2][7]= dspregs.W_Q2_0_0_7;
assign dspif.weight_bias[2][8]= dspregs.W_Q2_0_1_0;
assign dspif.weight_bias[2][9]= dspregs.W_Q2_0_1_1;
assign dspif.weight_bias[2][10]=dspregs.W_Q2_0_1_2;
assign dspif.weight_bias[2][11]=dspregs.W_Q2_0_1_3;
assign dspif.weight_bias[2][12]=dspregs.W_Q2_0_1_4;
assign dspif.weight_bias[2][13]=dspregs.W_Q2_0_1_5;
assign dspif.weight_bias[2][14]=dspregs.W_Q2_0_1_6;
assign dspif.weight_bias[2][15]=dspregs.W_Q2_0_1_7;
assign dspif.weight_bias[2][16]=dspregs.W_Q2_1_0_0;
assign dspif.weight_bias[2][17]=dspregs.W_Q2_1_0_1;
assign dspif.weight_bias[2][18]=dspregs.W_Q2_1_0_2;
assign dspif.weight_bias[2][19]=dspregs.W_Q2_1_0_3;
assign dspif.weight_bias[2][20]=dspregs.W_Q2_1_1_0;
assign dspif.weight_bias[2][21]=dspregs.W_Q2_1_1_1;
assign dspif.weight_bias[2][22]=dspregs.W_Q2_1_1_2;
assign dspif.weight_bias[2][23]=dspregs.W_Q2_1_1_3;
assign dspif.weight_bias[2][24]=dspregs.W_Q2_1_2_0;
assign dspif.weight_bias[2][25]=dspregs.W_Q2_1_2_1;
assign dspif.weight_bias[2][26]=dspregs.W_Q2_1_2_2;
assign dspif.weight_bias[2][27]=dspregs.W_Q2_1_2_3;
assign dspif.weight_bias[2][28]=dspregs.W_Q2_1_3_0;
assign dspif.weight_bias[2][29]=dspregs.W_Q2_1_3_1;
assign dspif.weight_bias[2][30]=dspregs.W_Q2_1_3_2;
assign dspif.weight_bias[2][31]=dspregs.W_Q2_1_3_3;
assign dspif.weight_bias[2][32]=dspregs.W_Q2_1_4_0;
assign dspif.weight_bias[2][33]=dspregs.W_Q2_1_4_1;
assign dspif.weight_bias[2][34]=dspregs.W_Q2_1_4_2;
assign dspif.weight_bias[2][35]=dspregs.W_Q2_1_4_3;
assign dspif.weight_bias[2][36]=dspregs.W_Q2_1_5_0;
assign dspif.weight_bias[2][37]=dspregs.W_Q2_1_5_1;
assign dspif.weight_bias[2][38]=dspregs.W_Q2_1_5_2;
assign dspif.weight_bias[2][39]=dspregs.W_Q2_1_5_3;
assign dspif.weight_bias[2][40]=dspregs.W_Q2_1_6_0;
assign dspif.weight_bias[2][41]=dspregs.W_Q2_1_6_1;
assign dspif.weight_bias[2][42]=dspregs.W_Q2_1_6_2;
assign dspif.weight_bias[2][43]=dspregs.W_Q2_1_6_3;
assign dspif.weight_bias[2][44]=dspregs.W_Q2_1_7_0;
assign dspif.weight_bias[2][45]=dspregs.W_Q2_1_7_1;
assign dspif.weight_bias[2][46]=dspregs.W_Q2_1_7_2;
assign dspif.weight_bias[2][47]=dspregs.W_Q2_1_7_3;
assign dspif.weight_bias[2][48]=dspregs.W_Q2_2_0_0;
assign dspif.weight_bias[2][49]=dspregs.W_Q2_2_1_0;
assign dspif.weight_bias[2][50]=dspregs.W_Q2_2_2_0;
assign dspif.weight_bias[2][51]=dspregs.W_Q2_2_3_0;
assign dspif.weight_bias[2][52]=dspregs.B_Q2_0_0;
assign dspif.weight_bias[2][53]=dspregs.B_Q2_0_1;
assign dspif.weight_bias[2][54]=dspregs.B_Q2_0_2;
assign dspif.weight_bias[2][55]=dspregs.B_Q2_0_3;
assign dspif.weight_bias[2][56]=dspregs.B_Q2_0_4;
assign dspif.weight_bias[2][57]=dspregs.B_Q2_0_5;
assign dspif.weight_bias[2][58]=dspregs.B_Q2_0_6;
assign dspif.weight_bias[2][59]=dspregs.B_Q2_0_7;
assign dspif.weight_bias[2][60]=dspregs.B_Q2_1_0;
assign dspif.weight_bias[2][61]=dspregs.B_Q2_1_1;
assign dspif.weight_bias[2][62]=dspregs.B_Q2_1_2;
assign dspif.weight_bias[2][63]=dspregs.B_Q2_1_3;
assign dspif.weight_bias[2][64]=dspregs.B_Q2_2_0;
assign dspif.weight_bias[3][0]= dspregs.W_Q3_0_0_0;
assign dspif.weight_bias[3][1]= dspregs.W_Q3_0_0_1;
assign dspif.weight_bias[3][2]= dspregs.W_Q3_0_0_2;
assign dspif.weight_bias[3][3]= dspregs.W_Q3_0_0_3;
assign dspif.weight_bias[3][4]= dspregs.W_Q3_0_0_4;
assign dspif.weight_bias[3][5]= dspregs.W_Q3_0_0_5;
assign dspif.weight_bias[3][6]= dspregs.W_Q3_0_0_6;
assign dspif.weight_bias[3][7]= dspregs.W_Q3_0_0_7;
assign dspif.weight_bias[3][8]= dspregs.W_Q3_0_1_0;
assign dspif.weight_bias[3][9]= dspregs.W_Q3_0_1_1;
assign dspif.weight_bias[3][10]=dspregs.W_Q3_0_1_2;
assign dspif.weight_bias[3][11]=dspregs.W_Q3_0_1_3;
assign dspif.weight_bias[3][12]=dspregs.W_Q3_0_1_4;
assign dspif.weight_bias[3][13]=dspregs.W_Q3_0_1_5;
assign dspif.weight_bias[3][14]=dspregs.W_Q3_0_1_6;
assign dspif.weight_bias[3][15]=dspregs.W_Q3_0_1_7;
assign dspif.weight_bias[3][16]=dspregs.W_Q3_1_0_0;
assign dspif.weight_bias[3][17]=dspregs.W_Q3_1_0_1;
assign dspif.weight_bias[3][18]=dspregs.W_Q3_1_0_2;
assign dspif.weight_bias[3][19]=dspregs.W_Q3_1_0_3;
assign dspif.weight_bias[3][20]=dspregs.W_Q3_1_1_0;
assign dspif.weight_bias[3][21]=dspregs.W_Q3_1_1_1;
assign dspif.weight_bias[3][22]=dspregs.W_Q3_1_1_2;
assign dspif.weight_bias[3][23]=dspregs.W_Q3_1_1_3;
assign dspif.weight_bias[3][24]=dspregs.W_Q3_1_2_0;
assign dspif.weight_bias[3][25]=dspregs.W_Q3_1_2_1;
assign dspif.weight_bias[3][26]=dspregs.W_Q3_1_2_2;
assign dspif.weight_bias[3][27]=dspregs.W_Q3_1_2_3;
assign dspif.weight_bias[3][28]=dspregs.W_Q3_1_3_0;
assign dspif.weight_bias[3][29]=dspregs.W_Q3_1_3_1;
assign dspif.weight_bias[3][30]=dspregs.W_Q3_1_3_2;
assign dspif.weight_bias[3][31]=dspregs.W_Q3_1_3_3;
assign dspif.weight_bias[3][32]=dspregs.W_Q3_1_4_0;
assign dspif.weight_bias[3][33]=dspregs.W_Q3_1_4_1;
assign dspif.weight_bias[3][34]=dspregs.W_Q3_1_4_2;
assign dspif.weight_bias[3][35]=dspregs.W_Q3_1_4_3;
assign dspif.weight_bias[3][36]=dspregs.W_Q3_1_5_0;
assign dspif.weight_bias[3][37]=dspregs.W_Q3_1_5_1;
assign dspif.weight_bias[3][38]=dspregs.W_Q3_1_5_2;
assign dspif.weight_bias[3][39]=dspregs.W_Q3_1_5_3;
assign dspif.weight_bias[3][40]=dspregs.W_Q3_1_6_0;
assign dspif.weight_bias[3][41]=dspregs.W_Q3_1_6_1;
assign dspif.weight_bias[3][42]=dspregs.W_Q3_1_6_2;
assign dspif.weight_bias[3][43]=dspregs.W_Q3_1_6_3;
assign dspif.weight_bias[3][44]=dspregs.W_Q3_1_7_0;
assign dspif.weight_bias[3][45]=dspregs.W_Q3_1_7_1;
assign dspif.weight_bias[3][46]=dspregs.W_Q3_1_7_2;
assign dspif.weight_bias[3][47]=dspregs.W_Q3_1_7_3;
assign dspif.weight_bias[3][48]=dspregs.W_Q3_2_0_0;
assign dspif.weight_bias[3][49]=dspregs.W_Q3_2_1_0;
assign dspif.weight_bias[3][50]=dspregs.W_Q3_2_2_0;
assign dspif.weight_bias[3][51]=dspregs.W_Q3_2_3_0;
assign dspif.weight_bias[3][52]=dspregs.B_Q3_0_0;
assign dspif.weight_bias[3][53]=dspregs.B_Q3_0_1;
assign dspif.weight_bias[3][54]=dspregs.B_Q3_0_2;
assign dspif.weight_bias[3][55]=dspregs.B_Q3_0_3;
assign dspif.weight_bias[3][56]=dspregs.B_Q3_0_4;
assign dspif.weight_bias[3][57]=dspregs.B_Q3_0_5;
assign dspif.weight_bias[3][58]=dspregs.B_Q3_0_6;
assign dspif.weight_bias[3][59]=dspregs.B_Q3_0_7;
assign dspif.weight_bias[3][60]=dspregs.B_Q3_1_0;
assign dspif.weight_bias[3][61]=dspregs.B_Q3_1_1;
assign dspif.weight_bias[3][62]=dspregs.B_Q3_1_2;
assign dspif.weight_bias[3][63]=dspregs.B_Q3_1_3;
assign dspif.weight_bias[3][64]=dspregs.B_Q3_2_0;
assign dspif.weight_bias[4][0]= dspregs.W_Q4_0_0_0;
assign dspif.weight_bias[4][1]= dspregs.W_Q4_0_0_1;
assign dspif.weight_bias[4][2]= dspregs.W_Q4_0_0_2;
assign dspif.weight_bias[4][3]= dspregs.W_Q4_0_0_3;
assign dspif.weight_bias[4][4]= dspregs.W_Q4_0_0_4;
assign dspif.weight_bias[4][5]= dspregs.W_Q4_0_0_5;
assign dspif.weight_bias[4][6]= dspregs.W_Q4_0_0_6;
assign dspif.weight_bias[4][7]= dspregs.W_Q4_0_0_7;
assign dspif.weight_bias[4][8]= dspregs.W_Q4_0_1_0;
assign dspif.weight_bias[4][9]= dspregs.W_Q4_0_1_1;
assign dspif.weight_bias[4][10]=dspregs.W_Q4_0_1_2;
assign dspif.weight_bias[4][11]=dspregs.W_Q4_0_1_3;
assign dspif.weight_bias[4][12]=dspregs.W_Q4_0_1_4;
assign dspif.weight_bias[4][13]=dspregs.W_Q4_0_1_5;
assign dspif.weight_bias[4][14]=dspregs.W_Q4_0_1_6;
assign dspif.weight_bias[4][15]=dspregs.W_Q4_0_1_7;
assign dspif.weight_bias[4][16]=dspregs.W_Q4_1_0_0;
assign dspif.weight_bias[4][17]=dspregs.W_Q4_1_0_1;
assign dspif.weight_bias[4][18]=dspregs.W_Q4_1_0_2;
assign dspif.weight_bias[4][19]=dspregs.W_Q4_1_0_3;
assign dspif.weight_bias[4][20]=dspregs.W_Q4_1_1_0;
assign dspif.weight_bias[4][21]=dspregs.W_Q4_1_1_1;
assign dspif.weight_bias[4][22]=dspregs.W_Q4_1_1_2;
assign dspif.weight_bias[4][23]=dspregs.W_Q4_1_1_3;
assign dspif.weight_bias[4][24]=dspregs.W_Q4_1_2_0;
assign dspif.weight_bias[4][25]=dspregs.W_Q4_1_2_1;
assign dspif.weight_bias[4][26]=dspregs.W_Q4_1_2_2;
assign dspif.weight_bias[4][27]=dspregs.W_Q4_1_2_3;
assign dspif.weight_bias[4][28]=dspregs.W_Q4_1_3_0;
assign dspif.weight_bias[4][29]=dspregs.W_Q4_1_3_1;
assign dspif.weight_bias[4][30]=dspregs.W_Q4_1_3_2;
assign dspif.weight_bias[4][31]=dspregs.W_Q4_1_3_3;
assign dspif.weight_bias[4][32]=dspregs.W_Q4_1_4_0;
assign dspif.weight_bias[4][33]=dspregs.W_Q4_1_4_1;
assign dspif.weight_bias[4][34]=dspregs.W_Q4_1_4_2;
assign dspif.weight_bias[4][35]=dspregs.W_Q4_1_4_3;
assign dspif.weight_bias[4][36]=dspregs.W_Q4_1_5_0;
assign dspif.weight_bias[4][37]=dspregs.W_Q4_1_5_1;
assign dspif.weight_bias[4][38]=dspregs.W_Q4_1_5_2;
assign dspif.weight_bias[4][39]=dspregs.W_Q4_1_5_3;
assign dspif.weight_bias[4][40]=dspregs.W_Q4_1_6_0;
assign dspif.weight_bias[4][41]=dspregs.W_Q4_1_6_1;
assign dspif.weight_bias[4][42]=dspregs.W_Q4_1_6_2;
assign dspif.weight_bias[4][43]=dspregs.W_Q4_1_6_3;
assign dspif.weight_bias[4][44]=dspregs.W_Q4_1_7_0;
assign dspif.weight_bias[4][45]=dspregs.W_Q4_1_7_1;
assign dspif.weight_bias[4][46]=dspregs.W_Q4_1_7_2;
assign dspif.weight_bias[4][47]=dspregs.W_Q4_1_7_3;
assign dspif.weight_bias[4][48]=dspregs.W_Q4_2_0_0;
assign dspif.weight_bias[4][49]=dspregs.W_Q4_2_1_0;
assign dspif.weight_bias[4][50]=dspregs.W_Q4_2_2_0;
assign dspif.weight_bias[4][51]=dspregs.W_Q4_2_3_0;
assign dspif.weight_bias[4][52]=dspregs.B_Q4_0_0;
assign dspif.weight_bias[4][53]=dspregs.B_Q4_0_1;
assign dspif.weight_bias[4][54]=dspregs.B_Q4_0_2;
assign dspif.weight_bias[4][55]=dspregs.B_Q4_0_3;
assign dspif.weight_bias[4][56]=dspregs.B_Q4_0_4;
assign dspif.weight_bias[4][57]=dspregs.B_Q4_0_5;
assign dspif.weight_bias[4][58]=dspregs.B_Q4_0_6;
assign dspif.weight_bias[4][59]=dspregs.B_Q4_0_7;
assign dspif.weight_bias[4][60]=dspregs.B_Q4_1_0;
assign dspif.weight_bias[4][61]=dspregs.B_Q4_1_1;
assign dspif.weight_bias[4][62]=dspregs.B_Q4_1_2;
assign dspif.weight_bias[4][63]=dspregs.B_Q4_1_3;
assign dspif.weight_bias[4][64]=dspregs.B_Q4_2_0;
assign dspif.weight_bias[5][0]= dspregs.W_Q5_0_0_0;
assign dspif.weight_bias[5][1]= dspregs.W_Q5_0_0_1;
assign dspif.weight_bias[5][2]= dspregs.W_Q5_0_0_2;
assign dspif.weight_bias[5][3]= dspregs.W_Q5_0_0_3;
assign dspif.weight_bias[5][4]= dspregs.W_Q5_0_0_4;
assign dspif.weight_bias[5][5]= dspregs.W_Q5_0_0_5;
assign dspif.weight_bias[5][6]= dspregs.W_Q5_0_0_6;
assign dspif.weight_bias[5][7]= dspregs.W_Q5_0_0_7;
assign dspif.weight_bias[5][8]= dspregs.W_Q5_0_1_0;
assign dspif.weight_bias[5][9]= dspregs.W_Q5_0_1_1;
assign dspif.weight_bias[5][10]=dspregs.W_Q5_0_1_2;
assign dspif.weight_bias[5][11]=dspregs.W_Q5_0_1_3;
assign dspif.weight_bias[5][12]=dspregs.W_Q5_0_1_4;
assign dspif.weight_bias[5][13]=dspregs.W_Q5_0_1_5;
assign dspif.weight_bias[5][14]=dspregs.W_Q5_0_1_6;
assign dspif.weight_bias[5][15]=dspregs.W_Q5_0_1_7;
assign dspif.weight_bias[5][16]=dspregs.W_Q5_1_0_0;
assign dspif.weight_bias[5][17]=dspregs.W_Q5_1_0_1;
assign dspif.weight_bias[5][18]=dspregs.W_Q5_1_0_2;
assign dspif.weight_bias[5][19]=dspregs.W_Q5_1_0_3;
assign dspif.weight_bias[5][20]=dspregs.W_Q5_1_1_0;
assign dspif.weight_bias[5][21]=dspregs.W_Q5_1_1_1;
assign dspif.weight_bias[5][22]=dspregs.W_Q5_1_1_2;
assign dspif.weight_bias[5][23]=dspregs.W_Q5_1_1_3;
assign dspif.weight_bias[5][24]=dspregs.W_Q5_1_2_0;
assign dspif.weight_bias[5][25]=dspregs.W_Q5_1_2_1;
assign dspif.weight_bias[5][26]=dspregs.W_Q5_1_2_2;
assign dspif.weight_bias[5][27]=dspregs.W_Q5_1_2_3;
assign dspif.weight_bias[5][28]=dspregs.W_Q5_1_3_0;
assign dspif.weight_bias[5][29]=dspregs.W_Q5_1_3_1;
assign dspif.weight_bias[5][30]=dspregs.W_Q5_1_3_2;
assign dspif.weight_bias[5][31]=dspregs.W_Q5_1_3_3;
assign dspif.weight_bias[5][32]=dspregs.W_Q5_1_4_0;
assign dspif.weight_bias[5][33]=dspregs.W_Q5_1_4_1;
assign dspif.weight_bias[5][34]=dspregs.W_Q5_1_4_2;
assign dspif.weight_bias[5][35]=dspregs.W_Q5_1_4_3;
assign dspif.weight_bias[5][36]=dspregs.W_Q5_1_5_0;
assign dspif.weight_bias[5][37]=dspregs.W_Q5_1_5_1;
assign dspif.weight_bias[5][38]=dspregs.W_Q5_1_5_2;
assign dspif.weight_bias[5][39]=dspregs.W_Q5_1_5_3;
assign dspif.weight_bias[5][40]=dspregs.W_Q5_1_6_0;
assign dspif.weight_bias[5][41]=dspregs.W_Q5_1_6_1;
assign dspif.weight_bias[5][42]=dspregs.W_Q5_1_6_2;
assign dspif.weight_bias[5][43]=dspregs.W_Q5_1_6_3;
assign dspif.weight_bias[5][44]=dspregs.W_Q5_1_7_0;
assign dspif.weight_bias[5][45]=dspregs.W_Q5_1_7_1;
assign dspif.weight_bias[5][46]=dspregs.W_Q5_1_7_2;
assign dspif.weight_bias[5][47]=dspregs.W_Q5_1_7_3;
assign dspif.weight_bias[5][48]=dspregs.W_Q5_2_0_0;
assign dspif.weight_bias[5][49]=dspregs.W_Q5_2_1_0;
assign dspif.weight_bias[5][50]=dspregs.W_Q5_2_2_0;
assign dspif.weight_bias[5][51]=dspregs.W_Q5_2_3_0;
assign dspif.weight_bias[5][52]=dspregs.B_Q5_0_0;
assign dspif.weight_bias[5][53]=dspregs.B_Q5_0_1;
assign dspif.weight_bias[5][54]=dspregs.B_Q5_0_2;
assign dspif.weight_bias[5][55]=dspregs.B_Q5_0_3;
assign dspif.weight_bias[5][56]=dspregs.B_Q5_0_4;
assign dspif.weight_bias[5][57]=dspregs.B_Q5_0_5;
assign dspif.weight_bias[5][58]=dspregs.B_Q5_0_6;
assign dspif.weight_bias[5][59]=dspregs.B_Q5_0_7;
assign dspif.weight_bias[5][60]=dspregs.B_Q5_1_0;
assign dspif.weight_bias[5][61]=dspregs.B_Q5_1_1;
assign dspif.weight_bias[5][62]=dspregs.B_Q5_1_2;
assign dspif.weight_bias[5][63]=dspregs.B_Q5_1_3;
assign dspif.weight_bias[5][64]=dspregs.B_Q5_2_0;
assign dspif.weight_bias[6][0]= dspregs.W_Q6_0_0_0;
assign dspif.weight_bias[6][1]= dspregs.W_Q6_0_0_1;
assign dspif.weight_bias[6][2]= dspregs.W_Q6_0_0_2;
assign dspif.weight_bias[6][3]= dspregs.W_Q6_0_0_3;
assign dspif.weight_bias[6][4]= dspregs.W_Q6_0_0_4;
assign dspif.weight_bias[6][5]= dspregs.W_Q6_0_0_5;
assign dspif.weight_bias[6][6]= dspregs.W_Q6_0_0_6;
assign dspif.weight_bias[6][7]= dspregs.W_Q6_0_0_7;
assign dspif.weight_bias[6][8]= dspregs.W_Q6_0_1_0;
assign dspif.weight_bias[6][9]= dspregs.W_Q6_0_1_1;
assign dspif.weight_bias[6][10]=dspregs.W_Q6_0_1_2;
assign dspif.weight_bias[6][11]=dspregs.W_Q6_0_1_3;
assign dspif.weight_bias[6][12]=dspregs.W_Q6_0_1_4;
assign dspif.weight_bias[6][13]=dspregs.W_Q6_0_1_5;
assign dspif.weight_bias[6][14]=dspregs.W_Q6_0_1_6;
assign dspif.weight_bias[6][15]=dspregs.W_Q6_0_1_7;
assign dspif.weight_bias[6][16]=dspregs.W_Q6_1_0_0;
assign dspif.weight_bias[6][17]=dspregs.W_Q6_1_0_1;
assign dspif.weight_bias[6][18]=dspregs.W_Q6_1_0_2;
assign dspif.weight_bias[6][19]=dspregs.W_Q6_1_0_3;
assign dspif.weight_bias[6][20]=dspregs.W_Q6_1_1_0;
assign dspif.weight_bias[6][21]=dspregs.W_Q6_1_1_1;
assign dspif.weight_bias[6][22]=dspregs.W_Q6_1_1_2;
assign dspif.weight_bias[6][23]=dspregs.W_Q6_1_1_3;
assign dspif.weight_bias[6][24]=dspregs.W_Q6_1_2_0;
assign dspif.weight_bias[6][25]=dspregs.W_Q6_1_2_1;
assign dspif.weight_bias[6][26]=dspregs.W_Q6_1_2_2;
assign dspif.weight_bias[6][27]=dspregs.W_Q6_1_2_3;
assign dspif.weight_bias[6][28]=dspregs.W_Q6_1_3_0;
assign dspif.weight_bias[6][29]=dspregs.W_Q6_1_3_1;
assign dspif.weight_bias[6][30]=dspregs.W_Q6_1_3_2;
assign dspif.weight_bias[6][31]=dspregs.W_Q6_1_3_3;
assign dspif.weight_bias[6][32]=dspregs.W_Q6_1_4_0;
assign dspif.weight_bias[6][33]=dspregs.W_Q6_1_4_1;
assign dspif.weight_bias[6][34]=dspregs.W_Q6_1_4_2;
assign dspif.weight_bias[6][35]=dspregs.W_Q6_1_4_3;
assign dspif.weight_bias[6][36]=dspregs.W_Q6_1_5_0;
assign dspif.weight_bias[6][37]=dspregs.W_Q6_1_5_1;
assign dspif.weight_bias[6][38]=dspregs.W_Q6_1_5_2;
assign dspif.weight_bias[6][39]=dspregs.W_Q6_1_5_3;
assign dspif.weight_bias[6][40]=dspregs.W_Q6_1_6_0;
assign dspif.weight_bias[6][41]=dspregs.W_Q6_1_6_1;
assign dspif.weight_bias[6][42]=dspregs.W_Q6_1_6_2;
assign dspif.weight_bias[6][43]=dspregs.W_Q6_1_6_3;
assign dspif.weight_bias[6][44]=dspregs.W_Q6_1_7_0;
assign dspif.weight_bias[6][45]=dspregs.W_Q6_1_7_1;
assign dspif.weight_bias[6][46]=dspregs.W_Q6_1_7_2;
assign dspif.weight_bias[6][47]=dspregs.W_Q6_1_7_3;
assign dspif.weight_bias[6][48]=dspregs.W_Q6_2_0_0;
assign dspif.weight_bias[6][49]=dspregs.W_Q6_2_1_0;
assign dspif.weight_bias[6][50]=dspregs.W_Q6_2_2_0;
assign dspif.weight_bias[6][51]=dspregs.W_Q6_2_3_0;
assign dspif.weight_bias[6][52]=dspregs.B_Q6_0_0;
assign dspif.weight_bias[6][53]=dspregs.B_Q6_0_1;
assign dspif.weight_bias[6][54]=dspregs.B_Q6_0_2;
assign dspif.weight_bias[6][55]=dspregs.B_Q6_0_3;
assign dspif.weight_bias[6][56]=dspregs.B_Q6_0_4;
assign dspif.weight_bias[6][57]=dspregs.B_Q6_0_5;
assign dspif.weight_bias[6][58]=dspregs.B_Q6_0_6;
assign dspif.weight_bias[6][59]=dspregs.B_Q6_0_7;
assign dspif.weight_bias[6][60]=dspregs.B_Q6_1_0;
assign dspif.weight_bias[6][61]=dspregs.B_Q6_1_1;
assign dspif.weight_bias[6][62]=dspregs.B_Q6_1_2;
assign dspif.weight_bias[6][63]=dspregs.B_Q6_1_3;
assign dspif.weight_bias[6][64]=dspregs.B_Q6_2_0;
assign dspif.weight_bias[7][0]= dspregs.W_Q7_0_0_0;
assign dspif.weight_bias[7][1]= dspregs.W_Q7_0_0_1;
assign dspif.weight_bias[7][2]= dspregs.W_Q7_0_0_2;
assign dspif.weight_bias[7][3]= dspregs.W_Q7_0_0_3;
assign dspif.weight_bias[7][4]= dspregs.W_Q7_0_0_4;
assign dspif.weight_bias[7][5]= dspregs.W_Q7_0_0_5;
assign dspif.weight_bias[7][6]= dspregs.W_Q7_0_0_6;
assign dspif.weight_bias[7][7]= dspregs.W_Q7_0_0_7;
assign dspif.weight_bias[7][8]= dspregs.W_Q7_0_1_0;
assign dspif.weight_bias[7][9]= dspregs.W_Q7_0_1_1;
assign dspif.weight_bias[7][10]=dspregs.W_Q7_0_1_2;
assign dspif.weight_bias[7][11]=dspregs.W_Q7_0_1_3;
assign dspif.weight_bias[7][12]=dspregs.W_Q7_0_1_4;
assign dspif.weight_bias[7][13]=dspregs.W_Q7_0_1_5;
assign dspif.weight_bias[7][14]=dspregs.W_Q7_0_1_6;
assign dspif.weight_bias[7][15]=dspregs.W_Q7_0_1_7;
assign dspif.weight_bias[7][16]=dspregs.W_Q7_1_0_0;
assign dspif.weight_bias[7][17]=dspregs.W_Q7_1_0_1;
assign dspif.weight_bias[7][18]=dspregs.W_Q7_1_0_2;
assign dspif.weight_bias[7][19]=dspregs.W_Q7_1_0_3;
assign dspif.weight_bias[7][20]=dspregs.W_Q7_1_1_0;
assign dspif.weight_bias[7][21]=dspregs.W_Q7_1_1_1;
assign dspif.weight_bias[7][22]=dspregs.W_Q7_1_1_2;
assign dspif.weight_bias[7][23]=dspregs.W_Q7_1_1_3;
assign dspif.weight_bias[7][24]=dspregs.W_Q7_1_2_0;
assign dspif.weight_bias[7][25]=dspregs.W_Q7_1_2_1;
assign dspif.weight_bias[7][26]=dspregs.W_Q7_1_2_2;
assign dspif.weight_bias[7][27]=dspregs.W_Q7_1_2_3;
assign dspif.weight_bias[7][28]=dspregs.W_Q7_1_3_0;
assign dspif.weight_bias[7][29]=dspregs.W_Q7_1_3_1;
assign dspif.weight_bias[7][30]=dspregs.W_Q7_1_3_2;
assign dspif.weight_bias[7][31]=dspregs.W_Q7_1_3_3;
assign dspif.weight_bias[7][32]=dspregs.W_Q7_1_4_0;
assign dspif.weight_bias[7][33]=dspregs.W_Q7_1_4_1;
assign dspif.weight_bias[7][34]=dspregs.W_Q7_1_4_2;
assign dspif.weight_bias[7][35]=dspregs.W_Q7_1_4_3;
assign dspif.weight_bias[7][36]=dspregs.W_Q7_1_5_0;
assign dspif.weight_bias[7][37]=dspregs.W_Q7_1_5_1;
assign dspif.weight_bias[7][38]=dspregs.W_Q7_1_5_2;
assign dspif.weight_bias[7][39]=dspregs.W_Q7_1_5_3;
assign dspif.weight_bias[7][40]=dspregs.W_Q7_1_6_0;
assign dspif.weight_bias[7][41]=dspregs.W_Q7_1_6_1;
assign dspif.weight_bias[7][42]=dspregs.W_Q7_1_6_2;
assign dspif.weight_bias[7][43]=dspregs.W_Q7_1_6_3;
assign dspif.weight_bias[7][44]=dspregs.W_Q7_1_7_0;
assign dspif.weight_bias[7][45]=dspregs.W_Q7_1_7_1;
assign dspif.weight_bias[7][46]=dspregs.W_Q7_1_7_2;
assign dspif.weight_bias[7][47]=dspregs.W_Q7_1_7_3;
assign dspif.weight_bias[7][48]=dspregs.W_Q7_2_0_0;
assign dspif.weight_bias[7][49]=dspregs.W_Q7_2_1_0;
assign dspif.weight_bias[7][50]=dspregs.W_Q7_2_2_0;
assign dspif.weight_bias[7][51]=dspregs.W_Q7_2_3_0;
assign dspif.weight_bias[7][52]=dspregs.B_Q7_0_0;
assign dspif.weight_bias[7][53]=dspregs.B_Q7_0_1;
assign dspif.weight_bias[7][54]=dspregs.B_Q7_0_2;
assign dspif.weight_bias[7][55]=dspregs.B_Q7_0_3;
assign dspif.weight_bias[7][56]=dspregs.B_Q7_0_4;
assign dspif.weight_bias[7][57]=dspregs.B_Q7_0_5;
assign dspif.weight_bias[7][58]=dspregs.B_Q7_0_6;
assign dspif.weight_bias[7][59]=dspregs.B_Q7_0_7;
assign dspif.weight_bias[7][60]=dspregs.B_Q7_1_0;
assign dspif.weight_bias[7][61]=dspregs.B_Q7_1_1;
assign dspif.weight_bias[7][62]=dspregs.B_Q7_1_2;
assign dspif.weight_bias[7][63]=dspregs.B_Q7_1_3;
assign dspif.weight_bias[7][64]=dspregs.B_Q7_2_0;

assign dspif.normalizer_min[0][0]=dspregs.min_Q0_I;
assign dspif.normalizer_min[0][1]=dspregs.min_Q0_Q;
assign dspif.normalizer_min[1][0]=dspregs.min_Q1_I;
assign dspif.normalizer_min[1][1]=dspregs.min_Q1_Q;
assign dspif.normalizer_min[2][0]=dspregs.min_Q2_I;
assign dspif.normalizer_min[2][1]=dspregs.min_Q2_Q;
assign dspif.normalizer_min[3][0]=dspregs.min_Q3_I;
assign dspif.normalizer_min[3][1]=dspregs.min_Q3_Q;
assign dspif.normalizer_min[4][0]=dspregs.min_Q4_I;
assign dspif.normalizer_min[4][1]=dspregs.min_Q4_Q;
assign dspif.normalizer_min[5][0]=dspregs.min_Q5_I;
assign dspif.normalizer_min[5][1]=dspregs.min_Q5_Q;
assign dspif.normalizer_min[6][0]=dspregs.min_Q6_I;
assign dspif.normalizer_min[6][1]=dspregs.min_Q6_Q;
assign dspif.normalizer_min[7][0]=dspregs.min_Q7_I;
assign dspif.normalizer_min[7][1]=dspregs.min_Q7_Q;
