.DAC00_M_AXIS_ACLK(DAC00_M_AXIS_ACLK)
    ,.DAC00_M_AXIS_ARESETN(DAC00_M_AXIS_ARESETN)
    ,.DAC00_M_AXIS_TREADY(DAC00_M_AXIS_TREADY)
    ,.DAC00_M_AXIS_TVALID(DAC00_M_AXIS_TVALID)
    ,.DAC00_M_AXIS_TDATA(DAC00_M_AXIS_TDATA)
    ,.DAC00_M_AXIS_TSTRB(DAC00_M_AXIS_TSTRB)
    ,.DAC00_M_AXIS_TLAST(DAC00_M_AXIS_TLAST)
,.clk_dac0(clk_dac0)
,.DAC01_M_AXIS_ACLK(DAC01_M_AXIS_ACLK)
    ,.DAC01_M_AXIS_ARESETN(DAC01_M_AXIS_ARESETN)
    ,.DAC01_M_AXIS_TREADY(DAC01_M_AXIS_TREADY)
    ,.DAC01_M_AXIS_TVALID(DAC01_M_AXIS_TVALID)
    ,.DAC01_M_AXIS_TDATA(DAC01_M_AXIS_TDATA)
    ,.DAC01_M_AXIS_TSTRB(DAC01_M_AXIS_TSTRB)
    ,.DAC01_M_AXIS_TLAST(DAC01_M_AXIS_TLAST)
,.DAC02_M_AXIS_ACLK(DAC02_M_AXIS_ACLK)
    ,.DAC02_M_AXIS_ARESETN(DAC02_M_AXIS_ARESETN)
    ,.DAC02_M_AXIS_TREADY(DAC02_M_AXIS_TREADY)
    ,.DAC02_M_AXIS_TVALID(DAC02_M_AXIS_TVALID)
    ,.DAC02_M_AXIS_TDATA(DAC02_M_AXIS_TDATA)
    ,.DAC02_M_AXIS_TSTRB(DAC02_M_AXIS_TSTRB)
    ,.DAC02_M_AXIS_TLAST(DAC02_M_AXIS_TLAST)
,.DAC03_M_AXIS_ACLK(DAC03_M_AXIS_ACLK)
    ,.DAC03_M_AXIS_ARESETN(DAC03_M_AXIS_ARESETN)
    ,.DAC03_M_AXIS_TREADY(DAC03_M_AXIS_TREADY)
    ,.DAC03_M_AXIS_TVALID(DAC03_M_AXIS_TVALID)
    ,.DAC03_M_AXIS_TDATA(DAC03_M_AXIS_TDATA)
    ,.DAC03_M_AXIS_TSTRB(DAC03_M_AXIS_TSTRB)
    ,.DAC03_M_AXIS_TLAST(DAC03_M_AXIS_TLAST)
,.DAC10_M_AXIS_ACLK(DAC10_M_AXIS_ACLK)
    ,.DAC10_M_AXIS_ARESETN(DAC10_M_AXIS_ARESETN)
    ,.DAC10_M_AXIS_TREADY(DAC10_M_AXIS_TREADY)
    ,.DAC10_M_AXIS_TVALID(DAC10_M_AXIS_TVALID)
    ,.DAC10_M_AXIS_TDATA(DAC10_M_AXIS_TDATA)
    ,.DAC10_M_AXIS_TSTRB(DAC10_M_AXIS_TSTRB)
    ,.DAC10_M_AXIS_TLAST(DAC10_M_AXIS_TLAST)
,.clk_dac1(clk_dac1)
,.DAC11_M_AXIS_ACLK(DAC11_M_AXIS_ACLK)
    ,.DAC11_M_AXIS_ARESETN(DAC11_M_AXIS_ARESETN)
    ,.DAC11_M_AXIS_TREADY(DAC11_M_AXIS_TREADY)
    ,.DAC11_M_AXIS_TVALID(DAC11_M_AXIS_TVALID)
    ,.DAC11_M_AXIS_TDATA(DAC11_M_AXIS_TDATA)
    ,.DAC11_M_AXIS_TSTRB(DAC11_M_AXIS_TSTRB)
    ,.DAC11_M_AXIS_TLAST(DAC11_M_AXIS_TLAST)
,.DAC12_M_AXIS_ACLK(DAC12_M_AXIS_ACLK)
    ,.DAC12_M_AXIS_ARESETN(DAC12_M_AXIS_ARESETN)
    ,.DAC12_M_AXIS_TREADY(DAC12_M_AXIS_TREADY)
    ,.DAC12_M_AXIS_TVALID(DAC12_M_AXIS_TVALID)
    ,.DAC12_M_AXIS_TDATA(DAC12_M_AXIS_TDATA)
    ,.DAC12_M_AXIS_TSTRB(DAC12_M_AXIS_TSTRB)
    ,.DAC12_M_AXIS_TLAST(DAC12_M_AXIS_TLAST)
,.DAC13_M_AXIS_ACLK(DAC13_M_AXIS_ACLK)
    ,.DAC13_M_AXIS_ARESETN(DAC13_M_AXIS_ARESETN)
    ,.DAC13_M_AXIS_TREADY(DAC13_M_AXIS_TREADY)
    ,.DAC13_M_AXIS_TVALID(DAC13_M_AXIS_TVALID)
    ,.DAC13_M_AXIS_TDATA(DAC13_M_AXIS_TDATA)
    ,.DAC13_M_AXIS_TSTRB(DAC13_M_AXIS_TSTRB)
    ,.DAC13_M_AXIS_TLAST(DAC13_M_AXIS_TLAST)
,.DAC20_M_AXIS_ACLK(DAC20_M_AXIS_ACLK)
    ,.DAC20_M_AXIS_ARESETN(DAC20_M_AXIS_ARESETN)
    ,.DAC20_M_AXIS_TREADY(DAC20_M_AXIS_TREADY)
    ,.DAC20_M_AXIS_TVALID(DAC20_M_AXIS_TVALID)
    ,.DAC20_M_AXIS_TDATA(DAC20_M_AXIS_TDATA)
    ,.DAC20_M_AXIS_TSTRB(DAC20_M_AXIS_TSTRB)
    ,.DAC20_M_AXIS_TLAST(DAC20_M_AXIS_TLAST)
,.clk_dac2(clk_dac2)
,.DAC21_M_AXIS_ACLK(DAC21_M_AXIS_ACLK)
    ,.DAC21_M_AXIS_ARESETN(DAC21_M_AXIS_ARESETN)
    ,.DAC21_M_AXIS_TREADY(DAC21_M_AXIS_TREADY)
    ,.DAC21_M_AXIS_TVALID(DAC21_M_AXIS_TVALID)
    ,.DAC21_M_AXIS_TDATA(DAC21_M_AXIS_TDATA)
    ,.DAC21_M_AXIS_TSTRB(DAC21_M_AXIS_TSTRB)
    ,.DAC21_M_AXIS_TLAST(DAC21_M_AXIS_TLAST)
,.DAC22_M_AXIS_ACLK(DAC22_M_AXIS_ACLK)
    ,.DAC22_M_AXIS_ARESETN(DAC22_M_AXIS_ARESETN)
    ,.DAC22_M_AXIS_TREADY(DAC22_M_AXIS_TREADY)
    ,.DAC22_M_AXIS_TVALID(DAC22_M_AXIS_TVALID)
    ,.DAC22_M_AXIS_TDATA(DAC22_M_AXIS_TDATA)
    ,.DAC22_M_AXIS_TSTRB(DAC22_M_AXIS_TSTRB)
    ,.DAC22_M_AXIS_TLAST(DAC22_M_AXIS_TLAST)
,.DAC23_M_AXIS_ACLK(DAC23_M_AXIS_ACLK)
    ,.DAC23_M_AXIS_ARESETN(DAC23_M_AXIS_ARESETN)
    ,.DAC23_M_AXIS_TREADY(DAC23_M_AXIS_TREADY)
    ,.DAC23_M_AXIS_TVALID(DAC23_M_AXIS_TVALID)
    ,.DAC23_M_AXIS_TDATA(DAC23_M_AXIS_TDATA)
    ,.DAC23_M_AXIS_TSTRB(DAC23_M_AXIS_TSTRB)
    ,.DAC23_M_AXIS_TLAST(DAC23_M_AXIS_TLAST)
,.DAC30_M_AXIS_ACLK(DAC30_M_AXIS_ACLK)
    ,.DAC30_M_AXIS_ARESETN(DAC30_M_AXIS_ARESETN)
    ,.DAC30_M_AXIS_TREADY(DAC30_M_AXIS_TREADY)
    ,.DAC30_M_AXIS_TVALID(DAC30_M_AXIS_TVALID)
    ,.DAC30_M_AXIS_TDATA(DAC30_M_AXIS_TDATA)
    ,.DAC30_M_AXIS_TSTRB(DAC30_M_AXIS_TSTRB)
    ,.DAC30_M_AXIS_TLAST(DAC30_M_AXIS_TLAST)
,.clk_dac3(clk_dac3)
,.DAC31_M_AXIS_ACLK(DAC31_M_AXIS_ACLK)
    ,.DAC31_M_AXIS_ARESETN(DAC31_M_AXIS_ARESETN)
    ,.DAC31_M_AXIS_TREADY(DAC31_M_AXIS_TREADY)
    ,.DAC31_M_AXIS_TVALID(DAC31_M_AXIS_TVALID)
    ,.DAC31_M_AXIS_TDATA(DAC31_M_AXIS_TDATA)
    ,.DAC31_M_AXIS_TSTRB(DAC31_M_AXIS_TSTRB)
    ,.DAC31_M_AXIS_TLAST(DAC31_M_AXIS_TLAST)
,.DAC32_M_AXIS_ACLK(DAC32_M_AXIS_ACLK)
    ,.DAC32_M_AXIS_ARESETN(DAC32_M_AXIS_ARESETN)
    ,.DAC32_M_AXIS_TREADY(DAC32_M_AXIS_TREADY)
    ,.DAC32_M_AXIS_TVALID(DAC32_M_AXIS_TVALID)
    ,.DAC32_M_AXIS_TDATA(DAC32_M_AXIS_TDATA)
    ,.DAC32_M_AXIS_TSTRB(DAC32_M_AXIS_TSTRB)
    ,.DAC32_M_AXIS_TLAST(DAC32_M_AXIS_TLAST)
,.DAC33_M_AXIS_ACLK(DAC33_M_AXIS_ACLK)
    ,.DAC33_M_AXIS_ARESETN(DAC33_M_AXIS_ARESETN)
    ,.DAC33_M_AXIS_TREADY(DAC33_M_AXIS_TREADY)
    ,.DAC33_M_AXIS_TVALID(DAC33_M_AXIS_TVALID)
    ,.DAC33_M_AXIS_TDATA(DAC33_M_AXIS_TDATA)
    ,.DAC33_M_AXIS_TSTRB(DAC33_M_AXIS_TSTRB)
    ,.DAC33_M_AXIS_TLAST(DAC33_M_AXIS_TLAST)
,.ADC00_S_AXIS_ACLK(ADC00_S_AXIS_ACLK)
    ,.ADC00_S_AXIS_ARESETN(ADC00_S_AXIS_ARESETN)
    ,.ADC00_S_AXIS_TREADY(ADC00_S_AXIS_TREADY)
    ,.ADC00_S_AXIS_TVALID(ADC00_S_AXIS_TVALID)
    ,.ADC00_S_AXIS_TDATA(ADC00_S_AXIS_TDATA)
    ,.ADC00_S_AXIS_TSTRB(ADC00_S_AXIS_TSTRB)
    ,.ADC00_S_AXIS_TLAST(ADC00_S_AXIS_TLAST)
,.clk_adc0(clk_adc0)
,.ADC01_S_AXIS_ACLK(ADC01_S_AXIS_ACLK)
    ,.ADC01_S_AXIS_ARESETN(ADC01_S_AXIS_ARESETN)
    ,.ADC01_S_AXIS_TREADY(ADC01_S_AXIS_TREADY)
    ,.ADC01_S_AXIS_TVALID(ADC01_S_AXIS_TVALID)
    ,.ADC01_S_AXIS_TDATA(ADC01_S_AXIS_TDATA)
    ,.ADC01_S_AXIS_TSTRB(ADC01_S_AXIS_TSTRB)
    ,.ADC01_S_AXIS_TLAST(ADC01_S_AXIS_TLAST)
,.ADC02_S_AXIS_ACLK(ADC02_S_AXIS_ACLK)
    ,.ADC02_S_AXIS_ARESETN(ADC02_S_AXIS_ARESETN)
    ,.ADC02_S_AXIS_TREADY(ADC02_S_AXIS_TREADY)
    ,.ADC02_S_AXIS_TVALID(ADC02_S_AXIS_TVALID)
    ,.ADC02_S_AXIS_TDATA(ADC02_S_AXIS_TDATA)
    ,.ADC02_S_AXIS_TSTRB(ADC02_S_AXIS_TSTRB)
    ,.ADC02_S_AXIS_TLAST(ADC02_S_AXIS_TLAST)
,.ADC03_S_AXIS_ACLK(ADC03_S_AXIS_ACLK)
    ,.ADC03_S_AXIS_ARESETN(ADC03_S_AXIS_ARESETN)
    ,.ADC03_S_AXIS_TREADY(ADC03_S_AXIS_TREADY)
    ,.ADC03_S_AXIS_TVALID(ADC03_S_AXIS_TVALID)
    ,.ADC03_S_AXIS_TDATA(ADC03_S_AXIS_TDATA)
    ,.ADC03_S_AXIS_TSTRB(ADC03_S_AXIS_TSTRB)
    ,.ADC03_S_AXIS_TLAST(ADC03_S_AXIS_TLAST)
,.ADC10_S_AXIS_ACLK(ADC10_S_AXIS_ACLK)
    ,.ADC10_S_AXIS_ARESETN(ADC10_S_AXIS_ARESETN)
    ,.ADC10_S_AXIS_TREADY(ADC10_S_AXIS_TREADY)
    ,.ADC10_S_AXIS_TVALID(ADC10_S_AXIS_TVALID)
    ,.ADC10_S_AXIS_TDATA(ADC10_S_AXIS_TDATA)
    ,.ADC10_S_AXIS_TSTRB(ADC10_S_AXIS_TSTRB)
    ,.ADC10_S_AXIS_TLAST(ADC10_S_AXIS_TLAST)
,.clk_adc1(clk_adc1)
,.ADC11_S_AXIS_ACLK(ADC11_S_AXIS_ACLK)
    ,.ADC11_S_AXIS_ARESETN(ADC11_S_AXIS_ARESETN)
    ,.ADC11_S_AXIS_TREADY(ADC11_S_AXIS_TREADY)
    ,.ADC11_S_AXIS_TVALID(ADC11_S_AXIS_TVALID)
    ,.ADC11_S_AXIS_TDATA(ADC11_S_AXIS_TDATA)
    ,.ADC11_S_AXIS_TSTRB(ADC11_S_AXIS_TSTRB)
    ,.ADC11_S_AXIS_TLAST(ADC11_S_AXIS_TLAST)
,.ADC12_S_AXIS_ACLK(ADC12_S_AXIS_ACLK)
    ,.ADC12_S_AXIS_ARESETN(ADC12_S_AXIS_ARESETN)
    ,.ADC12_S_AXIS_TREADY(ADC12_S_AXIS_TREADY)
    ,.ADC12_S_AXIS_TVALID(ADC12_S_AXIS_TVALID)
    ,.ADC12_S_AXIS_TDATA(ADC12_S_AXIS_TDATA)
    ,.ADC12_S_AXIS_TSTRB(ADC12_S_AXIS_TSTRB)
    ,.ADC12_S_AXIS_TLAST(ADC12_S_AXIS_TLAST)
,.ADC13_S_AXIS_ACLK(ADC13_S_AXIS_ACLK)
    ,.ADC13_S_AXIS_ARESETN(ADC13_S_AXIS_ARESETN)
    ,.ADC13_S_AXIS_TREADY(ADC13_S_AXIS_TREADY)
    ,.ADC13_S_AXIS_TVALID(ADC13_S_AXIS_TVALID)
    ,.ADC13_S_AXIS_TDATA(ADC13_S_AXIS_TDATA)
    ,.ADC13_S_AXIS_TSTRB(ADC13_S_AXIS_TSTRB)
    ,.ADC13_S_AXIS_TLAST(ADC13_S_AXIS_TLAST)
,.ADC20_S_AXIS_ACLK(ADC20_S_AXIS_ACLK)
    ,.ADC20_S_AXIS_ARESETN(ADC20_S_AXIS_ARESETN)
    ,.ADC20_S_AXIS_TREADY(ADC20_S_AXIS_TREADY)
    ,.ADC20_S_AXIS_TVALID(ADC20_S_AXIS_TVALID)
    ,.ADC20_S_AXIS_TDATA(ADC20_S_AXIS_TDATA)
    ,.ADC20_S_AXIS_TSTRB(ADC20_S_AXIS_TSTRB)
    ,.ADC20_S_AXIS_TLAST(ADC20_S_AXIS_TLAST)
,.clk_adc2(clk_adc2)
,.ADC21_S_AXIS_ACLK(ADC21_S_AXIS_ACLK)
    ,.ADC21_S_AXIS_ARESETN(ADC21_S_AXIS_ARESETN)
    ,.ADC21_S_AXIS_TREADY(ADC21_S_AXIS_TREADY)
    ,.ADC21_S_AXIS_TVALID(ADC21_S_AXIS_TVALID)
    ,.ADC21_S_AXIS_TDATA(ADC21_S_AXIS_TDATA)
    ,.ADC21_S_AXIS_TSTRB(ADC21_S_AXIS_TSTRB)
    ,.ADC21_S_AXIS_TLAST(ADC21_S_AXIS_TLAST)
,.ADC22_S_AXIS_ACLK(ADC22_S_AXIS_ACLK)
    ,.ADC22_S_AXIS_ARESETN(ADC22_S_AXIS_ARESETN)
    ,.ADC22_S_AXIS_TREADY(ADC22_S_AXIS_TREADY)
    ,.ADC22_S_AXIS_TVALID(ADC22_S_AXIS_TVALID)
    ,.ADC22_S_AXIS_TDATA(ADC22_S_AXIS_TDATA)
    ,.ADC22_S_AXIS_TSTRB(ADC22_S_AXIS_TSTRB)
    ,.ADC22_S_AXIS_TLAST(ADC22_S_AXIS_TLAST)
,.ADC23_S_AXIS_ACLK(ADC23_S_AXIS_ACLK)
    ,.ADC23_S_AXIS_ARESETN(ADC23_S_AXIS_ARESETN)
    ,.ADC23_S_AXIS_TREADY(ADC23_S_AXIS_TREADY)
    ,.ADC23_S_AXIS_TVALID(ADC23_S_AXIS_TVALID)
    ,.ADC23_S_AXIS_TDATA(ADC23_S_AXIS_TDATA)
    ,.ADC23_S_AXIS_TSTRB(ADC23_S_AXIS_TSTRB)
    ,.ADC23_S_AXIS_TLAST(ADC23_S_AXIS_TLAST)
,.ADC30_S_AXIS_ACLK(ADC30_S_AXIS_ACLK)
    ,.ADC30_S_AXIS_ARESETN(ADC30_S_AXIS_ARESETN)
    ,.ADC30_S_AXIS_TREADY(ADC30_S_AXIS_TREADY)
    ,.ADC30_S_AXIS_TVALID(ADC30_S_AXIS_TVALID)
    ,.ADC30_S_AXIS_TDATA(ADC30_S_AXIS_TDATA)
    ,.ADC30_S_AXIS_TSTRB(ADC30_S_AXIS_TSTRB)
    ,.ADC30_S_AXIS_TLAST(ADC30_S_AXIS_TLAST)
,.clk_adc3(clk_adc3)
,.ADC31_S_AXIS_ACLK(ADC31_S_AXIS_ACLK)
    ,.ADC31_S_AXIS_ARESETN(ADC31_S_AXIS_ARESETN)
    ,.ADC31_S_AXIS_TREADY(ADC31_S_AXIS_TREADY)
    ,.ADC31_S_AXIS_TVALID(ADC31_S_AXIS_TVALID)
    ,.ADC31_S_AXIS_TDATA(ADC31_S_AXIS_TDATA)
    ,.ADC31_S_AXIS_TSTRB(ADC31_S_AXIS_TSTRB)
    ,.ADC31_S_AXIS_TLAST(ADC31_S_AXIS_TLAST)
,.ADC32_S_AXIS_ACLK(ADC32_S_AXIS_ACLK)
    ,.ADC32_S_AXIS_ARESETN(ADC32_S_AXIS_ARESETN)
    ,.ADC32_S_AXIS_TREADY(ADC32_S_AXIS_TREADY)
    ,.ADC32_S_AXIS_TVALID(ADC32_S_AXIS_TVALID)
    ,.ADC32_S_AXIS_TDATA(ADC32_S_AXIS_TDATA)
    ,.ADC32_S_AXIS_TSTRB(ADC32_S_AXIS_TSTRB)
    ,.ADC32_S_AXIS_TLAST(ADC32_S_AXIS_TLAST)
,.ADC33_S_AXIS_ACLK(ADC33_S_AXIS_ACLK)
    ,.ADC33_S_AXIS_ARESETN(ADC33_S_AXIS_ARESETN)
    ,.ADC33_S_AXIS_TREADY(ADC33_S_AXIS_TREADY)
    ,.ADC33_S_AXIS_TVALID(ADC33_S_AXIS_TVALID)
    ,.ADC33_S_AXIS_TDATA(ADC33_S_AXIS_TDATA)
    ,.ADC33_S_AXIS_TSTRB(ADC33_S_AXIS_TSTRB)
    ,.ADC33_S_AXIS_TLAST(ADC33_S_AXIS_TLAST)