.cfgresetn0(cfgresetn0)
,.cfgresetn1(cfgresetn1)
,.cfgresetn2(cfgresetn2)
,.cfgresetn3(cfgresetn3)
,.cfgresetn4(cfgresetn4)
,.cfgresetn5(cfgresetn5)
,.cfgresetn6(cfgresetn6)
,.cfgresetn7(cfgresetn7)
,.dspresetn0(dspresetn0)
,.dspresetn1(dspresetn1)
,.dspresetn2(dspresetn2)
,.dspresetn3(dspresetn3)
,.dspresetn4(dspresetn4)
,.dspresetn5(dspresetn5)
,.dspresetn6(dspresetn6)
,.dspresetn7(dspresetn7)
,.dspresetn8(dspresetn8)
,.dspresetn9(dspresetn9)
,.dspresetn10(dspresetn10)
,.dspresetn11(dspresetn11)
,.dspresetn12(dspresetn12)
,.dspresetn13(dspresetn13)
,.dspresetn14(dspresetn14)
,.dspresetn15(dspresetn15)
,.dspresetn16(dspresetn16)
,.dspresetn17(dspresetn17)
,.dspresetn18(dspresetn18)
,.dspresetn19(dspresetn19)
,.dspresetn20(dspresetn20)
,.dspresetn21(dspresetn21)
,.dspresetn22(dspresetn22)
,.dspresetn23(dspresetn23)
,.dspresetn24(dspresetn24)
,.dspresetn25(dspresetn25)
,.dspresetn26(dspresetn26)
,.dspresetn27(dspresetn27)
,.dspresetn28(dspresetn28)
,.dspresetn29(dspresetn29)
,.dspresetn30(dspresetn30)
,.dspresetn31(dspresetn31)
,.dspresetn32(dspresetn32)
,.dspresetn33(dspresetn33)
,.dspresetn34(dspresetn34)
,.dspresetn35(dspresetn35)
,.dspresetn36(dspresetn36)
,.dspresetn37(dspresetn37)
,.dspresetn38(dspresetn38)
,.dspresetn39(dspresetn39)
,.dspresetn40(dspresetn40)
,.dspresetn41(dspresetn41)
,.psresetn0(psresetn0)
,.psresetn1(psresetn1)
,.psresetn2(psresetn2)
,.adc3resetn0(adc3resetn0)