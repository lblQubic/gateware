.dac00axis(dac00axis.master)
,.dac01axis(dac01axis.master)
,.dac02axis(dac02axis.master)
,.dac03axis(dac03axis.master)
,.dac10axis(dac10axis.master)
,.dac11axis(dac11axis.master)
,.dac12axis(dac12axis.master)
,.dac13axis(dac13axis.master)
,.dac20axis(dac20axis.master)
,.dac21axis(dac21axis.master)
,.dac22axis(dac22axis.master)
,.dac23axis(dac23axis.master)
,.dac30axis(dac30axis.master)
,.dac31axis(dac31axis.master)
,.dac32axis(dac32axis.master)
,.dac33axis(dac33axis.master)
,.adc00axis(adc00axis.slave)
,.adc01axis(adc01axis.slave)
,.adc02axis(adc02axis.slave)
,.adc03axis(adc03axis.slave)
,.adc10axis(adc10axis.slave)
,.adc11axis(adc11axis.slave)
,.adc12axis(adc12axis.slave)
,.adc13axis(adc13axis.slave)
,.adc20axis(adc20axis.slave)
,.adc21axis(adc21axis.slave)
,.adc22axis(adc22axis.slave)
,.adc23axis(adc23axis.slave)
,.adc30axis(adc30axis.slave)
,.adc31axis(adc31axis.slave)
,.adc32axis(adc32axis.slave)
,.adc33axis(adc33axis.slave)