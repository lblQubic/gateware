.INIT_acqbuf0(INIT_acqbuf0)
,.INIT_acqbuf1(INIT_acqbuf1)
,.INIT_command0(INIT_command0)
,.INIT_command1(INIT_command1)
,.INIT_command2(INIT_command2)
,.INIT_qdrvfreq0(INIT_qdrvfreq0)
,.INIT_qdrvfreq1(INIT_qdrvfreq1)
,.INIT_qdrvfreq2(INIT_qdrvfreq2)
,.INIT_rdrvfreq0(INIT_rdrvfreq0)
,.INIT_rdrvfreq1(INIT_rdrvfreq1)
,.INIT_rdrvfreq2(INIT_rdrvfreq2)
,.INIT_dacmon0(INIT_dacmon0)
,.INIT_dacmon1(INIT_dacmon1)
,.INIT_dacmon2(INIT_dacmon2)
,.INIT_dacmon3(INIT_dacmon3)
,.INIT_qdrvenv0(INIT_qdrvenv0)
,.INIT_qdrvenv1(INIT_qdrvenv1)
,.INIT_qdrvenv2(INIT_qdrvenv2)
,.INIT_rdloenv0(INIT_rdloenv0)
,.INIT_rdloenv1(INIT_rdloenv1)
,.INIT_rdloenv2(INIT_rdloenv2)
,.INIT_rdrvenv0(INIT_rdrvenv0)
,.INIT_rdrvenv1(INIT_rdrvenv1)
,.INIT_rdrvenv2(INIT_rdrvenv2)
,.INIT_accbuf0(INIT_accbuf0)
,.INIT_accbuf1(INIT_accbuf1)
,.INIT_accbuf2(INIT_accbuf2)
,.INIT_rdlofreq0(INIT_rdlofreq0)
,.INIT_rdlofreq1(INIT_rdlofreq1)
,.INIT_rdlofreq2(INIT_rdlofreq2)