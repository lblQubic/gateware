.ACCBUF0_clk(ACCBUF0_clk)
,.ACCBUF0_rst(ACCBUF0_rst)
,.ACCBUF0_addr(ACCBUF0_addr)
,.ACCBUF0_din(ACCBUF0_din)
,.ACCBUF0_dout(ACCBUF0_dout)
,.ACCBUF0_en(ACCBUF0_en)
,.ACCBUF0_we(ACCBUF0_we)

,.ACCBUF1_clk(ACCBUF1_clk)
,.ACCBUF1_rst(ACCBUF1_rst)
,.ACCBUF1_addr(ACCBUF1_addr)
,.ACCBUF1_din(ACCBUF1_din)
,.ACCBUF1_dout(ACCBUF1_dout)
,.ACCBUF1_en(ACCBUF1_en)
,.ACCBUF1_we(ACCBUF1_we)

,.ACCBUF2_clk(ACCBUF2_clk)
,.ACCBUF2_rst(ACCBUF2_rst)
,.ACCBUF2_addr(ACCBUF2_addr)
,.ACCBUF2_din(ACCBUF2_din)
,.ACCBUF2_dout(ACCBUF2_dout)
,.ACCBUF2_en(ACCBUF2_en)
,.ACCBUF2_we(ACCBUF2_we)

,.ACCBUF3_clk(ACCBUF3_clk)
,.ACCBUF3_rst(ACCBUF3_rst)
,.ACCBUF3_addr(ACCBUF3_addr)
,.ACCBUF3_din(ACCBUF3_din)
,.ACCBUF3_dout(ACCBUF3_dout)
,.ACCBUF3_en(ACCBUF3_en)
,.ACCBUF3_we(ACCBUF3_we)

,.ACCBUF4_clk(ACCBUF4_clk)
,.ACCBUF4_rst(ACCBUF4_rst)
,.ACCBUF4_addr(ACCBUF4_addr)
,.ACCBUF4_din(ACCBUF4_din)
,.ACCBUF4_dout(ACCBUF4_dout)
,.ACCBUF4_en(ACCBUF4_en)
,.ACCBUF4_we(ACCBUF4_we)

,.ACCBUF5_clk(ACCBUF5_clk)
,.ACCBUF5_rst(ACCBUF5_rst)
,.ACCBUF5_addr(ACCBUF5_addr)
,.ACCBUF5_din(ACCBUF5_din)
,.ACCBUF5_dout(ACCBUF5_dout)
,.ACCBUF5_en(ACCBUF5_en)
,.ACCBUF5_we(ACCBUF5_we)

,.ACCBUF6_clk(ACCBUF6_clk)
,.ACCBUF6_rst(ACCBUF6_rst)
,.ACCBUF6_addr(ACCBUF6_addr)
,.ACCBUF6_din(ACCBUF6_din)
,.ACCBUF6_dout(ACCBUF6_dout)
,.ACCBUF6_en(ACCBUF6_en)
,.ACCBUF6_we(ACCBUF6_we)

,.ACCBUF7_clk(ACCBUF7_clk)
,.ACCBUF7_rst(ACCBUF7_rst)
,.ACCBUF7_addr(ACCBUF7_addr)
,.ACCBUF7_din(ACCBUF7_din)
,.ACCBUF7_dout(ACCBUF7_dout)
,.ACCBUF7_en(ACCBUF7_en)
,.ACCBUF7_we(ACCBUF7_we)

,.ACQBUF0_clk(ACQBUF0_clk)
,.ACQBUF0_rst(ACQBUF0_rst)
,.ACQBUF0_addr(ACQBUF0_addr)
,.ACQBUF0_din(ACQBUF0_din)
,.ACQBUF0_dout(ACQBUF0_dout)
,.ACQBUF0_en(ACQBUF0_en)
,.ACQBUF0_we(ACQBUF0_we)

,.ACQBUF1_clk(ACQBUF1_clk)
,.ACQBUF1_rst(ACQBUF1_rst)
,.ACQBUF1_addr(ACQBUF1_addr)
,.ACQBUF1_din(ACQBUF1_din)
,.ACQBUF1_dout(ACQBUF1_dout)
,.ACQBUF1_en(ACQBUF1_en)
,.ACQBUF1_we(ACQBUF1_we)

,.COMMAND0_clk(COMMAND0_clk)
,.COMMAND0_rst(COMMAND0_rst)
,.COMMAND0_addr(COMMAND0_addr)
,.COMMAND0_din(COMMAND0_din)
,.COMMAND0_dout(COMMAND0_dout)
,.COMMAND0_en(COMMAND0_en)
,.COMMAND0_we(COMMAND0_we)

,.COMMAND1_clk(COMMAND1_clk)
,.COMMAND1_rst(COMMAND1_rst)
,.COMMAND1_addr(COMMAND1_addr)
,.COMMAND1_din(COMMAND1_din)
,.COMMAND1_dout(COMMAND1_dout)
,.COMMAND1_en(COMMAND1_en)
,.COMMAND1_we(COMMAND1_we)

,.COMMAND2_clk(COMMAND2_clk)
,.COMMAND2_rst(COMMAND2_rst)
,.COMMAND2_addr(COMMAND2_addr)
,.COMMAND2_din(COMMAND2_din)
,.COMMAND2_dout(COMMAND2_dout)
,.COMMAND2_en(COMMAND2_en)
,.COMMAND2_we(COMMAND2_we)

,.COMMAND3_clk(COMMAND3_clk)
,.COMMAND3_rst(COMMAND3_rst)
,.COMMAND3_addr(COMMAND3_addr)
,.COMMAND3_din(COMMAND3_din)
,.COMMAND3_dout(COMMAND3_dout)
,.COMMAND3_en(COMMAND3_en)
,.COMMAND3_we(COMMAND3_we)

,.COMMAND4_clk(COMMAND4_clk)
,.COMMAND4_rst(COMMAND4_rst)
,.COMMAND4_addr(COMMAND4_addr)
,.COMMAND4_din(COMMAND4_din)
,.COMMAND4_dout(COMMAND4_dout)
,.COMMAND4_en(COMMAND4_en)
,.COMMAND4_we(COMMAND4_we)

,.COMMAND5_clk(COMMAND5_clk)
,.COMMAND5_rst(COMMAND5_rst)
,.COMMAND5_addr(COMMAND5_addr)
,.COMMAND5_din(COMMAND5_din)
,.COMMAND5_dout(COMMAND5_dout)
,.COMMAND5_en(COMMAND5_en)
,.COMMAND5_we(COMMAND5_we)

,.COMMAND6_clk(COMMAND6_clk)
,.COMMAND6_rst(COMMAND6_rst)
,.COMMAND6_addr(COMMAND6_addr)
,.COMMAND6_din(COMMAND6_din)
,.COMMAND6_dout(COMMAND6_dout)
,.COMMAND6_en(COMMAND6_en)
,.COMMAND6_we(COMMAND6_we)

,.COMMAND7_clk(COMMAND7_clk)
,.COMMAND7_rst(COMMAND7_rst)
,.COMMAND7_addr(COMMAND7_addr)
,.COMMAND7_din(COMMAND7_din)
,.COMMAND7_dout(COMMAND7_dout)
,.COMMAND7_en(COMMAND7_en)
,.COMMAND7_we(COMMAND7_we)

,.DACMON0_clk(DACMON0_clk)
,.DACMON0_rst(DACMON0_rst)
,.DACMON0_addr(DACMON0_addr)
,.DACMON0_din(DACMON0_din)
,.DACMON0_dout(DACMON0_dout)
,.DACMON0_en(DACMON0_en)
,.DACMON0_we(DACMON0_we)

,.DACMON1_clk(DACMON1_clk)
,.DACMON1_rst(DACMON1_rst)
,.DACMON1_addr(DACMON1_addr)
,.DACMON1_din(DACMON1_din)
,.DACMON1_dout(DACMON1_dout)
,.DACMON1_en(DACMON1_en)
,.DACMON1_we(DACMON1_we)

,.DACMON2_clk(DACMON2_clk)
,.DACMON2_rst(DACMON2_rst)
,.DACMON2_addr(DACMON2_addr)
,.DACMON2_din(DACMON2_din)
,.DACMON2_dout(DACMON2_dout)
,.DACMON2_en(DACMON2_en)
,.DACMON2_we(DACMON2_we)

,.DACMON3_clk(DACMON3_clk)
,.DACMON3_rst(DACMON3_rst)
,.DACMON3_addr(DACMON3_addr)
,.DACMON3_din(DACMON3_din)
,.DACMON3_dout(DACMON3_dout)
,.DACMON3_en(DACMON3_en)
,.DACMON3_we(DACMON3_we)

,.QDRVENV0_clk(QDRVENV0_clk)
,.QDRVENV0_rst(QDRVENV0_rst)
,.QDRVENV0_addr(QDRVENV0_addr)
,.QDRVENV0_din(QDRVENV0_din)
,.QDRVENV0_dout(QDRVENV0_dout)
,.QDRVENV0_en(QDRVENV0_en)
,.QDRVENV0_we(QDRVENV0_we)

,.QDRVENV1_clk(QDRVENV1_clk)
,.QDRVENV1_rst(QDRVENV1_rst)
,.QDRVENV1_addr(QDRVENV1_addr)
,.QDRVENV1_din(QDRVENV1_din)
,.QDRVENV1_dout(QDRVENV1_dout)
,.QDRVENV1_en(QDRVENV1_en)
,.QDRVENV1_we(QDRVENV1_we)

,.QDRVENV2_clk(QDRVENV2_clk)
,.QDRVENV2_rst(QDRVENV2_rst)
,.QDRVENV2_addr(QDRVENV2_addr)
,.QDRVENV2_din(QDRVENV2_din)
,.QDRVENV2_dout(QDRVENV2_dout)
,.QDRVENV2_en(QDRVENV2_en)
,.QDRVENV2_we(QDRVENV2_we)

,.QDRVENV3_clk(QDRVENV3_clk)
,.QDRVENV3_rst(QDRVENV3_rst)
,.QDRVENV3_addr(QDRVENV3_addr)
,.QDRVENV3_din(QDRVENV3_din)
,.QDRVENV3_dout(QDRVENV3_dout)
,.QDRVENV3_en(QDRVENV3_en)
,.QDRVENV3_we(QDRVENV3_we)

,.QDRVENV4_clk(QDRVENV4_clk)
,.QDRVENV4_rst(QDRVENV4_rst)
,.QDRVENV4_addr(QDRVENV4_addr)
,.QDRVENV4_din(QDRVENV4_din)
,.QDRVENV4_dout(QDRVENV4_dout)
,.QDRVENV4_en(QDRVENV4_en)
,.QDRVENV4_we(QDRVENV4_we)

,.QDRVENV5_clk(QDRVENV5_clk)
,.QDRVENV5_rst(QDRVENV5_rst)
,.QDRVENV5_addr(QDRVENV5_addr)
,.QDRVENV5_din(QDRVENV5_din)
,.QDRVENV5_dout(QDRVENV5_dout)
,.QDRVENV5_en(QDRVENV5_en)
,.QDRVENV5_we(QDRVENV5_we)

,.QDRVENV6_clk(QDRVENV6_clk)
,.QDRVENV6_rst(QDRVENV6_rst)
,.QDRVENV6_addr(QDRVENV6_addr)
,.QDRVENV6_din(QDRVENV6_din)
,.QDRVENV6_dout(QDRVENV6_dout)
,.QDRVENV6_en(QDRVENV6_en)
,.QDRVENV6_we(QDRVENV6_we)

,.QDRVENV7_clk(QDRVENV7_clk)
,.QDRVENV7_rst(QDRVENV7_rst)
,.QDRVENV7_addr(QDRVENV7_addr)
,.QDRVENV7_din(QDRVENV7_din)
,.QDRVENV7_dout(QDRVENV7_dout)
,.QDRVENV7_en(QDRVENV7_en)
,.QDRVENV7_we(QDRVENV7_we)

,.QDRVFREQ0_clk(QDRVFREQ0_clk)
,.QDRVFREQ0_rst(QDRVFREQ0_rst)
,.QDRVFREQ0_addr(QDRVFREQ0_addr)
,.QDRVFREQ0_din(QDRVFREQ0_din)
,.QDRVFREQ0_dout(QDRVFREQ0_dout)
,.QDRVFREQ0_en(QDRVFREQ0_en)
,.QDRVFREQ0_we(QDRVFREQ0_we)

,.QDRVFREQ1_clk(QDRVFREQ1_clk)
,.QDRVFREQ1_rst(QDRVFREQ1_rst)
,.QDRVFREQ1_addr(QDRVFREQ1_addr)
,.QDRVFREQ1_din(QDRVFREQ1_din)
,.QDRVFREQ1_dout(QDRVFREQ1_dout)
,.QDRVFREQ1_en(QDRVFREQ1_en)
,.QDRVFREQ1_we(QDRVFREQ1_we)

,.QDRVFREQ2_clk(QDRVFREQ2_clk)
,.QDRVFREQ2_rst(QDRVFREQ2_rst)
,.QDRVFREQ2_addr(QDRVFREQ2_addr)
,.QDRVFREQ2_din(QDRVFREQ2_din)
,.QDRVFREQ2_dout(QDRVFREQ2_dout)
,.QDRVFREQ2_en(QDRVFREQ2_en)
,.QDRVFREQ2_we(QDRVFREQ2_we)

,.QDRVFREQ3_clk(QDRVFREQ3_clk)
,.QDRVFREQ3_rst(QDRVFREQ3_rst)
,.QDRVFREQ3_addr(QDRVFREQ3_addr)
,.QDRVFREQ3_din(QDRVFREQ3_din)
,.QDRVFREQ3_dout(QDRVFREQ3_dout)
,.QDRVFREQ3_en(QDRVFREQ3_en)
,.QDRVFREQ3_we(QDRVFREQ3_we)

,.QDRVFREQ4_clk(QDRVFREQ4_clk)
,.QDRVFREQ4_rst(QDRVFREQ4_rst)
,.QDRVFREQ4_addr(QDRVFREQ4_addr)
,.QDRVFREQ4_din(QDRVFREQ4_din)
,.QDRVFREQ4_dout(QDRVFREQ4_dout)
,.QDRVFREQ4_en(QDRVFREQ4_en)
,.QDRVFREQ4_we(QDRVFREQ4_we)

,.QDRVFREQ5_clk(QDRVFREQ5_clk)
,.QDRVFREQ5_rst(QDRVFREQ5_rst)
,.QDRVFREQ5_addr(QDRVFREQ5_addr)
,.QDRVFREQ5_din(QDRVFREQ5_din)
,.QDRVFREQ5_dout(QDRVFREQ5_dout)
,.QDRVFREQ5_en(QDRVFREQ5_en)
,.QDRVFREQ5_we(QDRVFREQ5_we)

,.QDRVFREQ6_clk(QDRVFREQ6_clk)
,.QDRVFREQ6_rst(QDRVFREQ6_rst)
,.QDRVFREQ6_addr(QDRVFREQ6_addr)
,.QDRVFREQ6_din(QDRVFREQ6_din)
,.QDRVFREQ6_dout(QDRVFREQ6_dout)
,.QDRVFREQ6_en(QDRVFREQ6_en)
,.QDRVFREQ6_we(QDRVFREQ6_we)

,.QDRVFREQ7_clk(QDRVFREQ7_clk)
,.QDRVFREQ7_rst(QDRVFREQ7_rst)
,.QDRVFREQ7_addr(QDRVFREQ7_addr)
,.QDRVFREQ7_din(QDRVFREQ7_din)
,.QDRVFREQ7_dout(QDRVFREQ7_dout)
,.QDRVFREQ7_en(QDRVFREQ7_en)
,.QDRVFREQ7_we(QDRVFREQ7_we)

,.RDLOENV0_clk(RDLOENV0_clk)
,.RDLOENV0_rst(RDLOENV0_rst)
,.RDLOENV0_addr(RDLOENV0_addr)
,.RDLOENV0_din(RDLOENV0_din)
,.RDLOENV0_dout(RDLOENV0_dout)
,.RDLOENV0_en(RDLOENV0_en)
,.RDLOENV0_we(RDLOENV0_we)

,.RDLOENV1_clk(RDLOENV1_clk)
,.RDLOENV1_rst(RDLOENV1_rst)
,.RDLOENV1_addr(RDLOENV1_addr)
,.RDLOENV1_din(RDLOENV1_din)
,.RDLOENV1_dout(RDLOENV1_dout)
,.RDLOENV1_en(RDLOENV1_en)
,.RDLOENV1_we(RDLOENV1_we)

,.RDLOENV2_clk(RDLOENV2_clk)
,.RDLOENV2_rst(RDLOENV2_rst)
,.RDLOENV2_addr(RDLOENV2_addr)
,.RDLOENV2_din(RDLOENV2_din)
,.RDLOENV2_dout(RDLOENV2_dout)
,.RDLOENV2_en(RDLOENV2_en)
,.RDLOENV2_we(RDLOENV2_we)

,.RDLOENV3_clk(RDLOENV3_clk)
,.RDLOENV3_rst(RDLOENV3_rst)
,.RDLOENV3_addr(RDLOENV3_addr)
,.RDLOENV3_din(RDLOENV3_din)
,.RDLOENV3_dout(RDLOENV3_dout)
,.RDLOENV3_en(RDLOENV3_en)
,.RDLOENV3_we(RDLOENV3_we)

,.RDLOENV4_clk(RDLOENV4_clk)
,.RDLOENV4_rst(RDLOENV4_rst)
,.RDLOENV4_addr(RDLOENV4_addr)
,.RDLOENV4_din(RDLOENV4_din)
,.RDLOENV4_dout(RDLOENV4_dout)
,.RDLOENV4_en(RDLOENV4_en)
,.RDLOENV4_we(RDLOENV4_we)

,.RDLOENV5_clk(RDLOENV5_clk)
,.RDLOENV5_rst(RDLOENV5_rst)
,.RDLOENV5_addr(RDLOENV5_addr)
,.RDLOENV5_din(RDLOENV5_din)
,.RDLOENV5_dout(RDLOENV5_dout)
,.RDLOENV5_en(RDLOENV5_en)
,.RDLOENV5_we(RDLOENV5_we)

,.RDLOENV6_clk(RDLOENV6_clk)
,.RDLOENV6_rst(RDLOENV6_rst)
,.RDLOENV6_addr(RDLOENV6_addr)
,.RDLOENV6_din(RDLOENV6_din)
,.RDLOENV6_dout(RDLOENV6_dout)
,.RDLOENV6_en(RDLOENV6_en)
,.RDLOENV6_we(RDLOENV6_we)

,.RDLOENV7_clk(RDLOENV7_clk)
,.RDLOENV7_rst(RDLOENV7_rst)
,.RDLOENV7_addr(RDLOENV7_addr)
,.RDLOENV7_din(RDLOENV7_din)
,.RDLOENV7_dout(RDLOENV7_dout)
,.RDLOENV7_en(RDLOENV7_en)
,.RDLOENV7_we(RDLOENV7_we)

,.RDLOFREQ0_clk(RDLOFREQ0_clk)
,.RDLOFREQ0_rst(RDLOFREQ0_rst)
,.RDLOFREQ0_addr(RDLOFREQ0_addr)
,.RDLOFREQ0_din(RDLOFREQ0_din)
,.RDLOFREQ0_dout(RDLOFREQ0_dout)
,.RDLOFREQ0_en(RDLOFREQ0_en)
,.RDLOFREQ0_we(RDLOFREQ0_we)

,.RDLOFREQ1_clk(RDLOFREQ1_clk)
,.RDLOFREQ1_rst(RDLOFREQ1_rst)
,.RDLOFREQ1_addr(RDLOFREQ1_addr)
,.RDLOFREQ1_din(RDLOFREQ1_din)
,.RDLOFREQ1_dout(RDLOFREQ1_dout)
,.RDLOFREQ1_en(RDLOFREQ1_en)
,.RDLOFREQ1_we(RDLOFREQ1_we)

,.RDLOFREQ2_clk(RDLOFREQ2_clk)
,.RDLOFREQ2_rst(RDLOFREQ2_rst)
,.RDLOFREQ2_addr(RDLOFREQ2_addr)
,.RDLOFREQ2_din(RDLOFREQ2_din)
,.RDLOFREQ2_dout(RDLOFREQ2_dout)
,.RDLOFREQ2_en(RDLOFREQ2_en)
,.RDLOFREQ2_we(RDLOFREQ2_we)

,.RDLOFREQ3_clk(RDLOFREQ3_clk)
,.RDLOFREQ3_rst(RDLOFREQ3_rst)
,.RDLOFREQ3_addr(RDLOFREQ3_addr)
,.RDLOFREQ3_din(RDLOFREQ3_din)
,.RDLOFREQ3_dout(RDLOFREQ3_dout)
,.RDLOFREQ3_en(RDLOFREQ3_en)
,.RDLOFREQ3_we(RDLOFREQ3_we)

,.RDLOFREQ4_clk(RDLOFREQ4_clk)
,.RDLOFREQ4_rst(RDLOFREQ4_rst)
,.RDLOFREQ4_addr(RDLOFREQ4_addr)
,.RDLOFREQ4_din(RDLOFREQ4_din)
,.RDLOFREQ4_dout(RDLOFREQ4_dout)
,.RDLOFREQ4_en(RDLOFREQ4_en)
,.RDLOFREQ4_we(RDLOFREQ4_we)

,.RDLOFREQ5_clk(RDLOFREQ5_clk)
,.RDLOFREQ5_rst(RDLOFREQ5_rst)
,.RDLOFREQ5_addr(RDLOFREQ5_addr)
,.RDLOFREQ5_din(RDLOFREQ5_din)
,.RDLOFREQ5_dout(RDLOFREQ5_dout)
,.RDLOFREQ5_en(RDLOFREQ5_en)
,.RDLOFREQ5_we(RDLOFREQ5_we)

,.RDLOFREQ6_clk(RDLOFREQ6_clk)
,.RDLOFREQ6_rst(RDLOFREQ6_rst)
,.RDLOFREQ6_addr(RDLOFREQ6_addr)
,.RDLOFREQ6_din(RDLOFREQ6_din)
,.RDLOFREQ6_dout(RDLOFREQ6_dout)
,.RDLOFREQ6_en(RDLOFREQ6_en)
,.RDLOFREQ6_we(RDLOFREQ6_we)

,.RDLOFREQ7_clk(RDLOFREQ7_clk)
,.RDLOFREQ7_rst(RDLOFREQ7_rst)
,.RDLOFREQ7_addr(RDLOFREQ7_addr)
,.RDLOFREQ7_din(RDLOFREQ7_din)
,.RDLOFREQ7_dout(RDLOFREQ7_dout)
,.RDLOFREQ7_en(RDLOFREQ7_en)
,.RDLOFREQ7_we(RDLOFREQ7_we)

,.RDRVENV0_clk(RDRVENV0_clk)
,.RDRVENV0_rst(RDRVENV0_rst)
,.RDRVENV0_addr(RDRVENV0_addr)
,.RDRVENV0_din(RDRVENV0_din)
,.RDRVENV0_dout(RDRVENV0_dout)
,.RDRVENV0_en(RDRVENV0_en)
,.RDRVENV0_we(RDRVENV0_we)

,.RDRVENV1_clk(RDRVENV1_clk)
,.RDRVENV1_rst(RDRVENV1_rst)
,.RDRVENV1_addr(RDRVENV1_addr)
,.RDRVENV1_din(RDRVENV1_din)
,.RDRVENV1_dout(RDRVENV1_dout)
,.RDRVENV1_en(RDRVENV1_en)
,.RDRVENV1_we(RDRVENV1_we)

,.RDRVENV2_clk(RDRVENV2_clk)
,.RDRVENV2_rst(RDRVENV2_rst)
,.RDRVENV2_addr(RDRVENV2_addr)
,.RDRVENV2_din(RDRVENV2_din)
,.RDRVENV2_dout(RDRVENV2_dout)
,.RDRVENV2_en(RDRVENV2_en)
,.RDRVENV2_we(RDRVENV2_we)

,.RDRVENV3_clk(RDRVENV3_clk)
,.RDRVENV3_rst(RDRVENV3_rst)
,.RDRVENV3_addr(RDRVENV3_addr)
,.RDRVENV3_din(RDRVENV3_din)
,.RDRVENV3_dout(RDRVENV3_dout)
,.RDRVENV3_en(RDRVENV3_en)
,.RDRVENV3_we(RDRVENV3_we)

,.RDRVENV4_clk(RDRVENV4_clk)
,.RDRVENV4_rst(RDRVENV4_rst)
,.RDRVENV4_addr(RDRVENV4_addr)
,.RDRVENV4_din(RDRVENV4_din)
,.RDRVENV4_dout(RDRVENV4_dout)
,.RDRVENV4_en(RDRVENV4_en)
,.RDRVENV4_we(RDRVENV4_we)

,.RDRVENV5_clk(RDRVENV5_clk)
,.RDRVENV5_rst(RDRVENV5_rst)
,.RDRVENV5_addr(RDRVENV5_addr)
,.RDRVENV5_din(RDRVENV5_din)
,.RDRVENV5_dout(RDRVENV5_dout)
,.RDRVENV5_en(RDRVENV5_en)
,.RDRVENV5_we(RDRVENV5_we)

,.RDRVENV6_clk(RDRVENV6_clk)
,.RDRVENV6_rst(RDRVENV6_rst)
,.RDRVENV6_addr(RDRVENV6_addr)
,.RDRVENV6_din(RDRVENV6_din)
,.RDRVENV6_dout(RDRVENV6_dout)
,.RDRVENV6_en(RDRVENV6_en)
,.RDRVENV6_we(RDRVENV6_we)

,.RDRVENV7_clk(RDRVENV7_clk)
,.RDRVENV7_rst(RDRVENV7_rst)
,.RDRVENV7_addr(RDRVENV7_addr)
,.RDRVENV7_din(RDRVENV7_din)
,.RDRVENV7_dout(RDRVENV7_dout)
,.RDRVENV7_en(RDRVENV7_en)
,.RDRVENV7_we(RDRVENV7_we)

,.RDRVFREQ0_clk(RDRVFREQ0_clk)
,.RDRVFREQ0_rst(RDRVFREQ0_rst)
,.RDRVFREQ0_addr(RDRVFREQ0_addr)
,.RDRVFREQ0_din(RDRVFREQ0_din)
,.RDRVFREQ0_dout(RDRVFREQ0_dout)
,.RDRVFREQ0_en(RDRVFREQ0_en)
,.RDRVFREQ0_we(RDRVFREQ0_we)

,.RDRVFREQ1_clk(RDRVFREQ1_clk)
,.RDRVFREQ1_rst(RDRVFREQ1_rst)
,.RDRVFREQ1_addr(RDRVFREQ1_addr)
,.RDRVFREQ1_din(RDRVFREQ1_din)
,.RDRVFREQ1_dout(RDRVFREQ1_dout)
,.RDRVFREQ1_en(RDRVFREQ1_en)
,.RDRVFREQ1_we(RDRVFREQ1_we)

,.RDRVFREQ2_clk(RDRVFREQ2_clk)
,.RDRVFREQ2_rst(RDRVFREQ2_rst)
,.RDRVFREQ2_addr(RDRVFREQ2_addr)
,.RDRVFREQ2_din(RDRVFREQ2_din)
,.RDRVFREQ2_dout(RDRVFREQ2_dout)
,.RDRVFREQ2_en(RDRVFREQ2_en)
,.RDRVFREQ2_we(RDRVFREQ2_we)

,.RDRVFREQ3_clk(RDRVFREQ3_clk)
,.RDRVFREQ3_rst(RDRVFREQ3_rst)
,.RDRVFREQ3_addr(RDRVFREQ3_addr)
,.RDRVFREQ3_din(RDRVFREQ3_din)
,.RDRVFREQ3_dout(RDRVFREQ3_dout)
,.RDRVFREQ3_en(RDRVFREQ3_en)
,.RDRVFREQ3_we(RDRVFREQ3_we)

,.RDRVFREQ4_clk(RDRVFREQ4_clk)
,.RDRVFREQ4_rst(RDRVFREQ4_rst)
,.RDRVFREQ4_addr(RDRVFREQ4_addr)
,.RDRVFREQ4_din(RDRVFREQ4_din)
,.RDRVFREQ4_dout(RDRVFREQ4_dout)
,.RDRVFREQ4_en(RDRVFREQ4_en)
,.RDRVFREQ4_we(RDRVFREQ4_we)

,.RDRVFREQ5_clk(RDRVFREQ5_clk)
,.RDRVFREQ5_rst(RDRVFREQ5_rst)
,.RDRVFREQ5_addr(RDRVFREQ5_addr)
,.RDRVFREQ5_din(RDRVFREQ5_din)
,.RDRVFREQ5_dout(RDRVFREQ5_dout)
,.RDRVFREQ5_en(RDRVFREQ5_en)
,.RDRVFREQ5_we(RDRVFREQ5_we)

,.RDRVFREQ6_clk(RDRVFREQ6_clk)
,.RDRVFREQ6_rst(RDRVFREQ6_rst)
,.RDRVFREQ6_addr(RDRVFREQ6_addr)
,.RDRVFREQ6_din(RDRVFREQ6_din)
,.RDRVFREQ6_dout(RDRVFREQ6_dout)
,.RDRVFREQ6_en(RDRVFREQ6_en)
,.RDRVFREQ6_we(RDRVFREQ6_we)

,.RDRVFREQ7_clk(RDRVFREQ7_clk)
,.RDRVFREQ7_rst(RDRVFREQ7_rst)
,.RDRVFREQ7_addr(RDRVFREQ7_addr)
,.RDRVFREQ7_din(RDRVFREQ7_din)
,.RDRVFREQ7_dout(RDRVFREQ7_dout)
,.RDRVFREQ7_en(RDRVFREQ7_en)
,.RDRVFREQ7_we(RDRVFREQ7_we)

,.SDBUF0_clk(SDBUF0_clk)
,.SDBUF0_rst(SDBUF0_rst)
,.SDBUF0_addr(SDBUF0_addr)
,.SDBUF0_din(SDBUF0_din)
,.SDBUF0_dout(SDBUF0_dout)
,.SDBUF0_en(SDBUF0_en)
,.SDBUF0_we(SDBUF0_we)

,.SDBUF1_clk(SDBUF1_clk)
,.SDBUF1_rst(SDBUF1_rst)
,.SDBUF1_addr(SDBUF1_addr)
,.SDBUF1_din(SDBUF1_din)
,.SDBUF1_dout(SDBUF1_dout)
,.SDBUF1_en(SDBUF1_en)
,.SDBUF1_we(SDBUF1_we)

,.SDBUF2_clk(SDBUF2_clk)
,.SDBUF2_rst(SDBUF2_rst)
,.SDBUF2_addr(SDBUF2_addr)
,.SDBUF2_din(SDBUF2_din)
,.SDBUF2_dout(SDBUF2_dout)
,.SDBUF2_en(SDBUF2_en)
,.SDBUF2_we(SDBUF2_we)

,.SDBUF3_clk(SDBUF3_clk)
,.SDBUF3_rst(SDBUF3_rst)
,.SDBUF3_addr(SDBUF3_addr)
,.SDBUF3_din(SDBUF3_din)
,.SDBUF3_dout(SDBUF3_dout)
,.SDBUF3_en(SDBUF3_en)
,.SDBUF3_we(SDBUF3_we)

,.SDBUF4_clk(SDBUF4_clk)
,.SDBUF4_rst(SDBUF4_rst)
,.SDBUF4_addr(SDBUF4_addr)
,.SDBUF4_din(SDBUF4_din)
,.SDBUF4_dout(SDBUF4_dout)
,.SDBUF4_en(SDBUF4_en)
,.SDBUF4_we(SDBUF4_we)

,.SDBUF5_clk(SDBUF5_clk)
,.SDBUF5_rst(SDBUF5_rst)
,.SDBUF5_addr(SDBUF5_addr)
,.SDBUF5_din(SDBUF5_din)
,.SDBUF5_dout(SDBUF5_dout)
,.SDBUF5_en(SDBUF5_en)
,.SDBUF5_we(SDBUF5_we)

,.SDBUF6_clk(SDBUF6_clk)
,.SDBUF6_rst(SDBUF6_rst)
,.SDBUF6_addr(SDBUF6_addr)
,.SDBUF6_din(SDBUF6_din)
,.SDBUF6_dout(SDBUF6_dout)
,.SDBUF6_en(SDBUF6_en)
,.SDBUF6_we(SDBUF6_we)

,.SDBUF7_clk(SDBUF7_clk)
,.SDBUF7_rst(SDBUF7_rst)
,.SDBUF7_addr(SDBUF7_addr)
,.SDBUF7_din(SDBUF7_din)
,.SDBUF7_dout(SDBUF7_dout)
,.SDBUF7_en(SDBUF7_en)
,.SDBUF7_we(SDBUF7_we)
