.acqbuf0_W(acqbuf0_W)
,.acqbuf1_W(acqbuf1_W)
,.command0_R(command0_R)
,.command1_R(command1_R)
,.command2_R(command2_R)
,.qdrvfreq0_R(qdrvfreq0_R)
,.qdrvfreq1_R(qdrvfreq1_R)
,.qdrvfreq2_R(qdrvfreq2_R)
,.rdrvfreq0_R(rdrvfreq0_R)
,.rdrvfreq1_R(rdrvfreq1_R)
,.rdrvfreq2_R(rdrvfreq2_R)
,.dacmon0_W(dacmon0_W)
,.dacmon1_W(dacmon1_W)
,.dacmon2_W(dacmon2_W)
,.dacmon3_W(dacmon3_W)
,.qdrvenv0_R(qdrvenv0_R)
,.qdrvenv1_R(qdrvenv1_R)
,.qdrvenv2_R(qdrvenv2_R)
,.rdloenv0_R(rdloenv0_R)
,.rdloenv1_R(rdloenv1_R)
,.rdloenv2_R(rdloenv2_R)
,.rdrvenv0_R(rdrvenv0_R)
,.rdrvenv1_R(rdrvenv1_R)
,.rdrvenv2_R(rdrvenv2_R)
,.accbuf0_W(accbuf0_W)
,.accbuf1_W(accbuf1_W)
,.accbuf2_W(accbuf2_W)
,.rdlofreq0_R(rdlofreq0_R)
,.rdlofreq1_R(rdlofreq1_R)
,.rdlofreq2_R(rdlofreq2_R)