interface ifdspregs #(parameter integer DATA_WIDTH = 32,parameter integer ADDR_WIDTH=24, parameter integer READDELAY=1)(    iflocalbus.lb lb
);
modport regs(input resetacc,stb_resetacc,amp,stb_amp,bramsel,stb_bramsel,coef00,stb_coef00,coef01,stb_coef01,coef02,stb_coef02,coef03,stb_coef03,coef10,stb_coef10,coef11,stb_coef11,coef12,stb_coef12,coef13,stb_coef13,coef20,stb_coef20,coef21,stb_coef21,coef22,stb_coef22,coef23,stb_coef23,coef30,stb_coef30,coef31,stb_coef31,coef32,stb_coef32,coef33,stb_coef33,dacsel,stb_dacsel,dspreset,stb_dspreset,nshot,stb_nshot,qdrvfreqsel,stb_qdrvfreqsel,rdlofreqsel,stb_rdlofreqsel,rdrvfreqsel,stb_rdrvfreqsel,reset_bram_read,stb_reset_bram_read,start,stb_start,test,stb_test,acqbufreset,stb_acqbufreset,dacmonreset,stb_dacmonreset,decimator,stb_decimator,acqchansel0,stb_acqchansel0,acqchansel1,stb_acqchansel1,dacmonchansel0,stb_dacmonchansel0,dacmonchansel1,stb_dacmonchansel1,dacmonchansel2,stb_dacmonchansel2,dacmonchansel3,stb_dacmonchansel3,delayaftertrig,stb_delayaftertrig,mixbb1sel,stb_mixbb1sel,mixbb2sel,stb_mixbb2sel,shift,stb_shift,W_Q0_0_0_0,stb_W_Q0_0_0_0,W_Q0_0_0_1,stb_W_Q0_0_0_1,W_Q0_0_0_2,stb_W_Q0_0_0_2,W_Q0_0_0_3,stb_W_Q0_0_0_3,W_Q0_0_0_4,stb_W_Q0_0_0_4,W_Q0_0_0_5,stb_W_Q0_0_0_5,W_Q0_0_0_6,stb_W_Q0_0_0_6,W_Q0_0_0_7,stb_W_Q0_0_0_7,W_Q0_0_1_0,stb_W_Q0_0_1_0,W_Q0_0_1_1,stb_W_Q0_0_1_1,W_Q0_0_1_2,stb_W_Q0_0_1_2,W_Q0_0_1_3,stb_W_Q0_0_1_3,W_Q0_0_1_4,stb_W_Q0_0_1_4,W_Q0_0_1_5,stb_W_Q0_0_1_5,W_Q0_0_1_6,stb_W_Q0_0_1_6,W_Q0_0_1_7,stb_W_Q0_0_1_7,W_Q0_1_0_0,stb_W_Q0_1_0_0,W_Q0_1_0_1,stb_W_Q0_1_0_1,W_Q0_1_0_2,stb_W_Q0_1_0_2,W_Q0_1_0_3,stb_W_Q0_1_0_3,W_Q0_1_1_0,stb_W_Q0_1_1_0,W_Q0_1_1_1,stb_W_Q0_1_1_1,W_Q0_1_1_2,stb_W_Q0_1_1_2,W_Q0_1_1_3,stb_W_Q0_1_1_3,W_Q0_1_2_0,stb_W_Q0_1_2_0,W_Q0_1_2_1,stb_W_Q0_1_2_1,W_Q0_1_2_2,stb_W_Q0_1_2_2,W_Q0_1_2_3,stb_W_Q0_1_2_3,W_Q0_1_3_0,stb_W_Q0_1_3_0,W_Q0_1_3_1,stb_W_Q0_1_3_1,W_Q0_1_3_2,stb_W_Q0_1_3_2,W_Q0_1_3_3,stb_W_Q0_1_3_3,W_Q0_1_4_0,stb_W_Q0_1_4_0,W_Q0_1_4_1,stb_W_Q0_1_4_1,W_Q0_1_4_2,stb_W_Q0_1_4_2,W_Q0_1_4_3,stb_W_Q0_1_4_3,W_Q0_1_5_0,stb_W_Q0_1_5_0,W_Q0_1_5_1,stb_W_Q0_1_5_1,W_Q0_1_5_2,stb_W_Q0_1_5_2,W_Q0_1_5_3,stb_W_Q0_1_5_3,W_Q0_1_6_0,stb_W_Q0_1_6_0,W_Q0_1_6_1,stb_W_Q0_1_6_1,W_Q0_1_6_2,stb_W_Q0_1_6_2,W_Q0_1_6_3,stb_W_Q0_1_6_3,W_Q0_1_7_0,stb_W_Q0_1_7_0,W_Q0_1_7_1,stb_W_Q0_1_7_1,W_Q0_1_7_2,stb_W_Q0_1_7_2,W_Q0_1_7_3,stb_W_Q0_1_7_3,W_Q0_2_0_0,stb_W_Q0_2_0_0,W_Q0_2_1_0,stb_W_Q0_2_1_0,W_Q0_2_2_0,stb_W_Q0_2_2_0,W_Q0_2_3_0,stb_W_Q0_2_3_0,B_Q0_0_0,stb_B_Q0_0_0,B_Q0_0_1,stb_B_Q0_0_1,B_Q0_0_2,stb_B_Q0_0_2,B_Q0_0_3,stb_B_Q0_0_3,B_Q0_0_4,stb_B_Q0_0_4,B_Q0_0_5,stb_B_Q0_0_5,B_Q0_0_6,stb_B_Q0_0_6,B_Q0_0_7,stb_B_Q0_0_7,B_Q0_1_0,stb_B_Q0_1_0,B_Q0_1_1,stb_B_Q0_1_1,B_Q0_1_2,stb_B_Q0_1_2,B_Q0_1_3,stb_B_Q0_1_3,B_Q0_2_0,stb_B_Q0_2_0,W_Q1_0_0_0,stb_W_Q1_0_0_0,W_Q1_0_0_1,stb_W_Q1_0_0_1,W_Q1_0_0_2,stb_W_Q1_0_0_2,W_Q1_0_0_3,stb_W_Q1_0_0_3,W_Q1_0_0_4,stb_W_Q1_0_0_4,W_Q1_0_0_5,stb_W_Q1_0_0_5,W_Q1_0_0_6,stb_W_Q1_0_0_6,W_Q1_0_0_7,stb_W_Q1_0_0_7,W_Q1_0_1_0,stb_W_Q1_0_1_0,W_Q1_0_1_1,stb_W_Q1_0_1_1,W_Q1_0_1_2,stb_W_Q1_0_1_2,W_Q1_0_1_3,stb_W_Q1_0_1_3,W_Q1_0_1_4,stb_W_Q1_0_1_4,W_Q1_0_1_5,stb_W_Q1_0_1_5,W_Q1_0_1_6,stb_W_Q1_0_1_6,W_Q1_0_1_7,stb_W_Q1_0_1_7,W_Q1_1_0_0,stb_W_Q1_1_0_0,W_Q1_1_0_1,stb_W_Q1_1_0_1,W_Q1_1_0_2,stb_W_Q1_1_0_2,W_Q1_1_0_3,stb_W_Q1_1_0_3,W_Q1_1_1_0,stb_W_Q1_1_1_0,W_Q1_1_1_1,stb_W_Q1_1_1_1,W_Q1_1_1_2,stb_W_Q1_1_1_2,W_Q1_1_1_3,stb_W_Q1_1_1_3,W_Q1_1_2_0,stb_W_Q1_1_2_0,W_Q1_1_2_1,stb_W_Q1_1_2_1,W_Q1_1_2_2,stb_W_Q1_1_2_2,W_Q1_1_2_3,stb_W_Q1_1_2_3,W_Q1_1_3_0,stb_W_Q1_1_3_0,W_Q1_1_3_1,stb_W_Q1_1_3_1,W_Q1_1_3_2,stb_W_Q1_1_3_2,W_Q1_1_3_3,stb_W_Q1_1_3_3,W_Q1_1_4_0,stb_W_Q1_1_4_0,W_Q1_1_4_1,stb_W_Q1_1_4_1,W_Q1_1_4_2,stb_W_Q1_1_4_2,W_Q1_1_4_3,stb_W_Q1_1_4_3,W_Q1_1_5_0,stb_W_Q1_1_5_0,W_Q1_1_5_1,stb_W_Q1_1_5_1,W_Q1_1_5_2,stb_W_Q1_1_5_2,W_Q1_1_5_3,stb_W_Q1_1_5_3,W_Q1_1_6_0,stb_W_Q1_1_6_0,W_Q1_1_6_1,stb_W_Q1_1_6_1,W_Q1_1_6_2,stb_W_Q1_1_6_2,W_Q1_1_6_3,stb_W_Q1_1_6_3,W_Q1_1_7_0,stb_W_Q1_1_7_0,W_Q1_1_7_1,stb_W_Q1_1_7_1,W_Q1_1_7_2,stb_W_Q1_1_7_2,W_Q1_1_7_3,stb_W_Q1_1_7_3,W_Q1_2_0_0,stb_W_Q1_2_0_0,W_Q1_2_1_0,stb_W_Q1_2_1_0,W_Q1_2_2_0,stb_W_Q1_2_2_0,W_Q1_2_3_0,stb_W_Q1_2_3_0,B_Q1_0_0,stb_B_Q1_0_0,B_Q1_0_1,stb_B_Q1_0_1,B_Q1_0_2,stb_B_Q1_0_2,B_Q1_0_3,stb_B_Q1_0_3,B_Q1_0_4,stb_B_Q1_0_4,B_Q1_0_5,stb_B_Q1_0_5,B_Q1_0_6,stb_B_Q1_0_6,B_Q1_0_7,stb_B_Q1_0_7,B_Q1_1_0,stb_B_Q1_1_0,B_Q1_1_1,stb_B_Q1_1_1,B_Q1_1_2,stb_B_Q1_1_2,B_Q1_1_3,stb_B_Q1_1_3,B_Q1_2_0,stb_B_Q1_2_0,W_Q2_0_0_0,stb_W_Q2_0_0_0,W_Q2_0_0_1,stb_W_Q2_0_0_1,W_Q2_0_0_2,stb_W_Q2_0_0_2,W_Q2_0_0_3,stb_W_Q2_0_0_3,W_Q2_0_0_4,stb_W_Q2_0_0_4,W_Q2_0_0_5,stb_W_Q2_0_0_5,W_Q2_0_0_6,stb_W_Q2_0_0_6,W_Q2_0_0_7,stb_W_Q2_0_0_7,W_Q2_0_1_0,stb_W_Q2_0_1_0,W_Q2_0_1_1,stb_W_Q2_0_1_1,W_Q2_0_1_2,stb_W_Q2_0_1_2,W_Q2_0_1_3,stb_W_Q2_0_1_3,W_Q2_0_1_4,stb_W_Q2_0_1_4,W_Q2_0_1_5,stb_W_Q2_0_1_5,W_Q2_0_1_6,stb_W_Q2_0_1_6,W_Q2_0_1_7,stb_W_Q2_0_1_7,W_Q2_1_0_0,stb_W_Q2_1_0_0,W_Q2_1_0_1,stb_W_Q2_1_0_1,W_Q2_1_0_2,stb_W_Q2_1_0_2,W_Q2_1_0_3,stb_W_Q2_1_0_3,W_Q2_1_1_0,stb_W_Q2_1_1_0,W_Q2_1_1_1,stb_W_Q2_1_1_1,W_Q2_1_1_2,stb_W_Q2_1_1_2,W_Q2_1_1_3,stb_W_Q2_1_1_3,W_Q2_1_2_0,stb_W_Q2_1_2_0,W_Q2_1_2_1,stb_W_Q2_1_2_1,W_Q2_1_2_2,stb_W_Q2_1_2_2,W_Q2_1_2_3,stb_W_Q2_1_2_3,W_Q2_1_3_0,stb_W_Q2_1_3_0,W_Q2_1_3_1,stb_W_Q2_1_3_1,W_Q2_1_3_2,stb_W_Q2_1_3_2,W_Q2_1_3_3,stb_W_Q2_1_3_3,W_Q2_1_4_0,stb_W_Q2_1_4_0,W_Q2_1_4_1,stb_W_Q2_1_4_1,W_Q2_1_4_2,stb_W_Q2_1_4_2,W_Q2_1_4_3,stb_W_Q2_1_4_3,W_Q2_1_5_0,stb_W_Q2_1_5_0,W_Q2_1_5_1,stb_W_Q2_1_5_1,W_Q2_1_5_2,stb_W_Q2_1_5_2,W_Q2_1_5_3,stb_W_Q2_1_5_3,W_Q2_1_6_0,stb_W_Q2_1_6_0,W_Q2_1_6_1,stb_W_Q2_1_6_1,W_Q2_1_6_2,stb_W_Q2_1_6_2,W_Q2_1_6_3,stb_W_Q2_1_6_3,W_Q2_1_7_0,stb_W_Q2_1_7_0,W_Q2_1_7_1,stb_W_Q2_1_7_1,W_Q2_1_7_2,stb_W_Q2_1_7_2,W_Q2_1_7_3,stb_W_Q2_1_7_3,W_Q2_2_0_0,stb_W_Q2_2_0_0,W_Q2_2_1_0,stb_W_Q2_2_1_0,W_Q2_2_2_0,stb_W_Q2_2_2_0,W_Q2_2_3_0,stb_W_Q2_2_3_0,B_Q2_0_0,stb_B_Q2_0_0,B_Q2_0_1,stb_B_Q2_0_1,B_Q2_0_2,stb_B_Q2_0_2,B_Q2_0_3,stb_B_Q2_0_3,B_Q2_0_4,stb_B_Q2_0_4,B_Q2_0_5,stb_B_Q2_0_5,B_Q2_0_6,stb_B_Q2_0_6,B_Q2_0_7,stb_B_Q2_0_7,B_Q2_1_0,stb_B_Q2_1_0,B_Q2_1_1,stb_B_Q2_1_1,B_Q2_1_2,stb_B_Q2_1_2,B_Q2_1_3,stb_B_Q2_1_3,B_Q2_2_0,stb_B_Q2_2_0,W_Q3_0_0_0,stb_W_Q3_0_0_0,W_Q3_0_0_1,stb_W_Q3_0_0_1,W_Q3_0_0_2,stb_W_Q3_0_0_2,W_Q3_0_0_3,stb_W_Q3_0_0_3,W_Q3_0_0_4,stb_W_Q3_0_0_4,W_Q3_0_0_5,stb_W_Q3_0_0_5,W_Q3_0_0_6,stb_W_Q3_0_0_6,W_Q3_0_0_7,stb_W_Q3_0_0_7,W_Q3_0_1_0,stb_W_Q3_0_1_0,W_Q3_0_1_1,stb_W_Q3_0_1_1,W_Q3_0_1_2,stb_W_Q3_0_1_2,W_Q3_0_1_3,stb_W_Q3_0_1_3,W_Q3_0_1_4,stb_W_Q3_0_1_4,W_Q3_0_1_5,stb_W_Q3_0_1_5,W_Q3_0_1_6,stb_W_Q3_0_1_6,W_Q3_0_1_7,stb_W_Q3_0_1_7,W_Q3_1_0_0,stb_W_Q3_1_0_0,W_Q3_1_0_1,stb_W_Q3_1_0_1,W_Q3_1_0_2,stb_W_Q3_1_0_2,W_Q3_1_0_3,stb_W_Q3_1_0_3,W_Q3_1_1_0,stb_W_Q3_1_1_0,W_Q3_1_1_1,stb_W_Q3_1_1_1,W_Q3_1_1_2,stb_W_Q3_1_1_2,W_Q3_1_1_3,stb_W_Q3_1_1_3,W_Q3_1_2_0,stb_W_Q3_1_2_0,W_Q3_1_2_1,stb_W_Q3_1_2_1,W_Q3_1_2_2,stb_W_Q3_1_2_2,W_Q3_1_2_3,stb_W_Q3_1_2_3,W_Q3_1_3_0,stb_W_Q3_1_3_0,W_Q3_1_3_1,stb_W_Q3_1_3_1,W_Q3_1_3_2,stb_W_Q3_1_3_2,W_Q3_1_3_3,stb_W_Q3_1_3_3,W_Q3_1_4_0,stb_W_Q3_1_4_0,W_Q3_1_4_1,stb_W_Q3_1_4_1,W_Q3_1_4_2,stb_W_Q3_1_4_2,W_Q3_1_4_3,stb_W_Q3_1_4_3,W_Q3_1_5_0,stb_W_Q3_1_5_0,W_Q3_1_5_1,stb_W_Q3_1_5_1,W_Q3_1_5_2,stb_W_Q3_1_5_2,W_Q3_1_5_3,stb_W_Q3_1_5_3,W_Q3_1_6_0,stb_W_Q3_1_6_0,W_Q3_1_6_1,stb_W_Q3_1_6_1,W_Q3_1_6_2,stb_W_Q3_1_6_2,W_Q3_1_6_3,stb_W_Q3_1_6_3,W_Q3_1_7_0,stb_W_Q3_1_7_0,W_Q3_1_7_1,stb_W_Q3_1_7_1,W_Q3_1_7_2,stb_W_Q3_1_7_2,W_Q3_1_7_3,stb_W_Q3_1_7_3,W_Q3_2_0_0,stb_W_Q3_2_0_0,W_Q3_2_1_0,stb_W_Q3_2_1_0,W_Q3_2_2_0,stb_W_Q3_2_2_0,W_Q3_2_3_0,stb_W_Q3_2_3_0,B_Q3_0_0,stb_B_Q3_0_0,B_Q3_0_1,stb_B_Q3_0_1,B_Q3_0_2,stb_B_Q3_0_2,B_Q3_0_3,stb_B_Q3_0_3,B_Q3_0_4,stb_B_Q3_0_4,B_Q3_0_5,stb_B_Q3_0_5,B_Q3_0_6,stb_B_Q3_0_6,B_Q3_0_7,stb_B_Q3_0_7,B_Q3_1_0,stb_B_Q3_1_0,B_Q3_1_1,stb_B_Q3_1_1,B_Q3_1_2,stb_B_Q3_1_2,B_Q3_1_3,stb_B_Q3_1_3,B_Q3_2_0,stb_B_Q3_2_0,W_Q4_0_0_0,stb_W_Q4_0_0_0,W_Q4_0_0_1,stb_W_Q4_0_0_1,W_Q4_0_0_2,stb_W_Q4_0_0_2,W_Q4_0_0_3,stb_W_Q4_0_0_3,W_Q4_0_0_4,stb_W_Q4_0_0_4,W_Q4_0_0_5,stb_W_Q4_0_0_5,W_Q4_0_0_6,stb_W_Q4_0_0_6,W_Q4_0_0_7,stb_W_Q4_0_0_7,W_Q4_0_1_0,stb_W_Q4_0_1_0,W_Q4_0_1_1,stb_W_Q4_0_1_1,W_Q4_0_1_2,stb_W_Q4_0_1_2,W_Q4_0_1_3,stb_W_Q4_0_1_3,W_Q4_0_1_4,stb_W_Q4_0_1_4,W_Q4_0_1_5,stb_W_Q4_0_1_5,W_Q4_0_1_6,stb_W_Q4_0_1_6,W_Q4_0_1_7,stb_W_Q4_0_1_7,W_Q4_1_0_0,stb_W_Q4_1_0_0,W_Q4_1_0_1,stb_W_Q4_1_0_1,W_Q4_1_0_2,stb_W_Q4_1_0_2,W_Q4_1_0_3,stb_W_Q4_1_0_3,W_Q4_1_1_0,stb_W_Q4_1_1_0,W_Q4_1_1_1,stb_W_Q4_1_1_1,W_Q4_1_1_2,stb_W_Q4_1_1_2,W_Q4_1_1_3,stb_W_Q4_1_1_3,W_Q4_1_2_0,stb_W_Q4_1_2_0,W_Q4_1_2_1,stb_W_Q4_1_2_1,W_Q4_1_2_2,stb_W_Q4_1_2_2,W_Q4_1_2_3,stb_W_Q4_1_2_3,W_Q4_1_3_0,stb_W_Q4_1_3_0,W_Q4_1_3_1,stb_W_Q4_1_3_1,W_Q4_1_3_2,stb_W_Q4_1_3_2,W_Q4_1_3_3,stb_W_Q4_1_3_3,W_Q4_1_4_0,stb_W_Q4_1_4_0,W_Q4_1_4_1,stb_W_Q4_1_4_1,W_Q4_1_4_2,stb_W_Q4_1_4_2,W_Q4_1_4_3,stb_W_Q4_1_4_3,W_Q4_1_5_0,stb_W_Q4_1_5_0,W_Q4_1_5_1,stb_W_Q4_1_5_1,W_Q4_1_5_2,stb_W_Q4_1_5_2,W_Q4_1_5_3,stb_W_Q4_1_5_3,W_Q4_1_6_0,stb_W_Q4_1_6_0,W_Q4_1_6_1,stb_W_Q4_1_6_1,W_Q4_1_6_2,stb_W_Q4_1_6_2,W_Q4_1_6_3,stb_W_Q4_1_6_3,W_Q4_1_7_0,stb_W_Q4_1_7_0,W_Q4_1_7_1,stb_W_Q4_1_7_1,W_Q4_1_7_2,stb_W_Q4_1_7_2,W_Q4_1_7_3,stb_W_Q4_1_7_3,W_Q4_2_0_0,stb_W_Q4_2_0_0,W_Q4_2_1_0,stb_W_Q4_2_1_0,W_Q4_2_2_0,stb_W_Q4_2_2_0,W_Q4_2_3_0,stb_W_Q4_2_3_0,B_Q4_0_0,stb_B_Q4_0_0,B_Q4_0_1,stb_B_Q4_0_1,B_Q4_0_2,stb_B_Q4_0_2,B_Q4_0_3,stb_B_Q4_0_3,B_Q4_0_4,stb_B_Q4_0_4,B_Q4_0_5,stb_B_Q4_0_5,B_Q4_0_6,stb_B_Q4_0_6,B_Q4_0_7,stb_B_Q4_0_7,B_Q4_1_0,stb_B_Q4_1_0,B_Q4_1_1,stb_B_Q4_1_1,B_Q4_1_2,stb_B_Q4_1_2,B_Q4_1_3,stb_B_Q4_1_3,B_Q4_2_0,stb_B_Q4_2_0,W_Q5_0_0_0,stb_W_Q5_0_0_0,W_Q5_0_0_1,stb_W_Q5_0_0_1,W_Q5_0_0_2,stb_W_Q5_0_0_2,W_Q5_0_0_3,stb_W_Q5_0_0_3,W_Q5_0_0_4,stb_W_Q5_0_0_4,W_Q5_0_0_5,stb_W_Q5_0_0_5,W_Q5_0_0_6,stb_W_Q5_0_0_6,W_Q5_0_0_7,stb_W_Q5_0_0_7,W_Q5_0_1_0,stb_W_Q5_0_1_0,W_Q5_0_1_1,stb_W_Q5_0_1_1,W_Q5_0_1_2,stb_W_Q5_0_1_2,W_Q5_0_1_3,stb_W_Q5_0_1_3,W_Q5_0_1_4,stb_W_Q5_0_1_4,W_Q5_0_1_5,stb_W_Q5_0_1_5,W_Q5_0_1_6,stb_W_Q5_0_1_6,W_Q5_0_1_7,stb_W_Q5_0_1_7,W_Q5_1_0_0,stb_W_Q5_1_0_0,W_Q5_1_0_1,stb_W_Q5_1_0_1,W_Q5_1_0_2,stb_W_Q5_1_0_2,W_Q5_1_0_3,stb_W_Q5_1_0_3,W_Q5_1_1_0,stb_W_Q5_1_1_0,W_Q5_1_1_1,stb_W_Q5_1_1_1,W_Q5_1_1_2,stb_W_Q5_1_1_2,W_Q5_1_1_3,stb_W_Q5_1_1_3,W_Q5_1_2_0,stb_W_Q5_1_2_0,W_Q5_1_2_1,stb_W_Q5_1_2_1,W_Q5_1_2_2,stb_W_Q5_1_2_2,W_Q5_1_2_3,stb_W_Q5_1_2_3,W_Q5_1_3_0,stb_W_Q5_1_3_0,W_Q5_1_3_1,stb_W_Q5_1_3_1,W_Q5_1_3_2,stb_W_Q5_1_3_2,W_Q5_1_3_3,stb_W_Q5_1_3_3,W_Q5_1_4_0,stb_W_Q5_1_4_0,W_Q5_1_4_1,stb_W_Q5_1_4_1,W_Q5_1_4_2,stb_W_Q5_1_4_2,W_Q5_1_4_3,stb_W_Q5_1_4_3,W_Q5_1_5_0,stb_W_Q5_1_5_0,W_Q5_1_5_1,stb_W_Q5_1_5_1,W_Q5_1_5_2,stb_W_Q5_1_5_2,W_Q5_1_5_3,stb_W_Q5_1_5_3,W_Q5_1_6_0,stb_W_Q5_1_6_0,W_Q5_1_6_1,stb_W_Q5_1_6_1,W_Q5_1_6_2,stb_W_Q5_1_6_2,W_Q5_1_6_3,stb_W_Q5_1_6_3,W_Q5_1_7_0,stb_W_Q5_1_7_0,W_Q5_1_7_1,stb_W_Q5_1_7_1,W_Q5_1_7_2,stb_W_Q5_1_7_2,W_Q5_1_7_3,stb_W_Q5_1_7_3,W_Q5_2_0_0,stb_W_Q5_2_0_0,W_Q5_2_1_0,stb_W_Q5_2_1_0,W_Q5_2_2_0,stb_W_Q5_2_2_0,W_Q5_2_3_0,stb_W_Q5_2_3_0,B_Q5_0_0,stb_B_Q5_0_0,B_Q5_0_1,stb_B_Q5_0_1,B_Q5_0_2,stb_B_Q5_0_2,B_Q5_0_3,stb_B_Q5_0_3,B_Q5_0_4,stb_B_Q5_0_4,B_Q5_0_5,stb_B_Q5_0_5,B_Q5_0_6,stb_B_Q5_0_6,B_Q5_0_7,stb_B_Q5_0_7,B_Q5_1_0,stb_B_Q5_1_0,B_Q5_1_1,stb_B_Q5_1_1,B_Q5_1_2,stb_B_Q5_1_2,B_Q5_1_3,stb_B_Q5_1_3,B_Q5_2_0,stb_B_Q5_2_0,W_Q6_0_0_0,stb_W_Q6_0_0_0,W_Q6_0_0_1,stb_W_Q6_0_0_1,W_Q6_0_0_2,stb_W_Q6_0_0_2,W_Q6_0_0_3,stb_W_Q6_0_0_3,W_Q6_0_0_4,stb_W_Q6_0_0_4,W_Q6_0_0_5,stb_W_Q6_0_0_5,W_Q6_0_0_6,stb_W_Q6_0_0_6,W_Q6_0_0_7,stb_W_Q6_0_0_7,W_Q6_0_1_0,stb_W_Q6_0_1_0,W_Q6_0_1_1,stb_W_Q6_0_1_1,W_Q6_0_1_2,stb_W_Q6_0_1_2,W_Q6_0_1_3,stb_W_Q6_0_1_3,W_Q6_0_1_4,stb_W_Q6_0_1_4,W_Q6_0_1_5,stb_W_Q6_0_1_5,W_Q6_0_1_6,stb_W_Q6_0_1_6,W_Q6_0_1_7,stb_W_Q6_0_1_7,W_Q6_1_0_0,stb_W_Q6_1_0_0,W_Q6_1_0_1,stb_W_Q6_1_0_1,W_Q6_1_0_2,stb_W_Q6_1_0_2,W_Q6_1_0_3,stb_W_Q6_1_0_3,W_Q6_1_1_0,stb_W_Q6_1_1_0,W_Q6_1_1_1,stb_W_Q6_1_1_1,W_Q6_1_1_2,stb_W_Q6_1_1_2,W_Q6_1_1_3,stb_W_Q6_1_1_3,W_Q6_1_2_0,stb_W_Q6_1_2_0,W_Q6_1_2_1,stb_W_Q6_1_2_1,W_Q6_1_2_2,stb_W_Q6_1_2_2,W_Q6_1_2_3,stb_W_Q6_1_2_3,W_Q6_1_3_0,stb_W_Q6_1_3_0,W_Q6_1_3_1,stb_W_Q6_1_3_1,W_Q6_1_3_2,stb_W_Q6_1_3_2,W_Q6_1_3_3,stb_W_Q6_1_3_3,W_Q6_1_4_0,stb_W_Q6_1_4_0,W_Q6_1_4_1,stb_W_Q6_1_4_1,W_Q6_1_4_2,stb_W_Q6_1_4_2,W_Q6_1_4_3,stb_W_Q6_1_4_3,W_Q6_1_5_0,stb_W_Q6_1_5_0,W_Q6_1_5_1,stb_W_Q6_1_5_1,W_Q6_1_5_2,stb_W_Q6_1_5_2,W_Q6_1_5_3,stb_W_Q6_1_5_3,W_Q6_1_6_0,stb_W_Q6_1_6_0,W_Q6_1_6_1,stb_W_Q6_1_6_1,W_Q6_1_6_2,stb_W_Q6_1_6_2,W_Q6_1_6_3,stb_W_Q6_1_6_3,W_Q6_1_7_0,stb_W_Q6_1_7_0,W_Q6_1_7_1,stb_W_Q6_1_7_1,W_Q6_1_7_2,stb_W_Q6_1_7_2,W_Q6_1_7_3,stb_W_Q6_1_7_3,W_Q6_2_0_0,stb_W_Q6_2_0_0,W_Q6_2_1_0,stb_W_Q6_2_1_0,W_Q6_2_2_0,stb_W_Q6_2_2_0,W_Q6_2_3_0,stb_W_Q6_2_3_0,B_Q6_0_0,stb_B_Q6_0_0,B_Q6_0_1,stb_B_Q6_0_1,B_Q6_0_2,stb_B_Q6_0_2,B_Q6_0_3,stb_B_Q6_0_3,B_Q6_0_4,stb_B_Q6_0_4,B_Q6_0_5,stb_B_Q6_0_5,B_Q6_0_6,stb_B_Q6_0_6,B_Q6_0_7,stb_B_Q6_0_7,B_Q6_1_0,stb_B_Q6_1_0,B_Q6_1_1,stb_B_Q6_1_1,B_Q6_1_2,stb_B_Q6_1_2,B_Q6_1_3,stb_B_Q6_1_3,B_Q6_2_0,stb_B_Q6_2_0,W_Q7_0_0_0,stb_W_Q7_0_0_0,W_Q7_0_0_1,stb_W_Q7_0_0_1,W_Q7_0_0_2,stb_W_Q7_0_0_2,W_Q7_0_0_3,stb_W_Q7_0_0_3,W_Q7_0_0_4,stb_W_Q7_0_0_4,W_Q7_0_0_5,stb_W_Q7_0_0_5,W_Q7_0_0_6,stb_W_Q7_0_0_6,W_Q7_0_0_7,stb_W_Q7_0_0_7,W_Q7_0_1_0,stb_W_Q7_0_1_0,W_Q7_0_1_1,stb_W_Q7_0_1_1,W_Q7_0_1_2,stb_W_Q7_0_1_2,W_Q7_0_1_3,stb_W_Q7_0_1_3,W_Q7_0_1_4,stb_W_Q7_0_1_4,W_Q7_0_1_5,stb_W_Q7_0_1_5,W_Q7_0_1_6,stb_W_Q7_0_1_6,W_Q7_0_1_7,stb_W_Q7_0_1_7,W_Q7_1_0_0,stb_W_Q7_1_0_0,W_Q7_1_0_1,stb_W_Q7_1_0_1,W_Q7_1_0_2,stb_W_Q7_1_0_2,W_Q7_1_0_3,stb_W_Q7_1_0_3,W_Q7_1_1_0,stb_W_Q7_1_1_0,W_Q7_1_1_1,stb_W_Q7_1_1_1,W_Q7_1_1_2,stb_W_Q7_1_1_2,W_Q7_1_1_3,stb_W_Q7_1_1_3,W_Q7_1_2_0,stb_W_Q7_1_2_0,W_Q7_1_2_1,stb_W_Q7_1_2_1,W_Q7_1_2_2,stb_W_Q7_1_2_2,W_Q7_1_2_3,stb_W_Q7_1_2_3,W_Q7_1_3_0,stb_W_Q7_1_3_0,W_Q7_1_3_1,stb_W_Q7_1_3_1,W_Q7_1_3_2,stb_W_Q7_1_3_2,W_Q7_1_3_3,stb_W_Q7_1_3_3,W_Q7_1_4_0,stb_W_Q7_1_4_0,W_Q7_1_4_1,stb_W_Q7_1_4_1,W_Q7_1_4_2,stb_W_Q7_1_4_2,W_Q7_1_4_3,stb_W_Q7_1_4_3,W_Q7_1_5_0,stb_W_Q7_1_5_0,W_Q7_1_5_1,stb_W_Q7_1_5_1,W_Q7_1_5_2,stb_W_Q7_1_5_2,W_Q7_1_5_3,stb_W_Q7_1_5_3,W_Q7_1_6_0,stb_W_Q7_1_6_0,W_Q7_1_6_1,stb_W_Q7_1_6_1,W_Q7_1_6_2,stb_W_Q7_1_6_2,W_Q7_1_6_3,stb_W_Q7_1_6_3,W_Q7_1_7_0,stb_W_Q7_1_7_0,W_Q7_1_7_1,stb_W_Q7_1_7_1,W_Q7_1_7_2,stb_W_Q7_1_7_2,W_Q7_1_7_3,stb_W_Q7_1_7_3,W_Q7_2_0_0,stb_W_Q7_2_0_0,W_Q7_2_1_0,stb_W_Q7_2_1_0,W_Q7_2_2_0,stb_W_Q7_2_2_0,W_Q7_2_3_0,stb_W_Q7_2_3_0,B_Q7_0_0,stb_B_Q7_0_0,B_Q7_0_1,stb_B_Q7_0_1,B_Q7_0_2,stb_B_Q7_0_2,B_Q7_0_3,stb_B_Q7_0_3,B_Q7_0_4,stb_B_Q7_0_4,B_Q7_0_5,stb_B_Q7_0_5,B_Q7_0_6,stb_B_Q7_0_6,B_Q7_0_7,stb_B_Q7_0_7,B_Q7_1_0,stb_B_Q7_1_0,B_Q7_1_1,stb_B_Q7_1_1,B_Q7_1_2,stb_B_Q7_1_2,B_Q7_1_3,stb_B_Q7_1_3,B_Q7_2_0,stb_B_Q7_2_0,min_Q0_I,stb_min_Q0_I,min_Q0_Q,stb_min_Q0_Q,min_Q1_I,stb_min_Q1_I,min_Q1_Q,stb_min_Q1_Q,min_Q2_I,stb_min_Q2_I,min_Q2_Q,stb_min_Q2_Q,min_Q3_I,stb_min_Q3_I,min_Q3_Q,stb_min_Q3_Q,min_Q4_I,stb_min_Q4_I,min_Q4_Q,stb_min_Q4_Q,min_Q5_I,stb_min_Q5_I,min_Q5_Q,stb_min_Q5_Q,min_Q6_I,stb_min_Q6_I,min_Q6_Q,stb_min_Q6_Q,min_Q7_I,stb_min_Q7_I,min_Q7_Q,stb_min_Q7_Q
,output addr_accbuf_mon0,addr_accbuf_mon1,addr_accbuf_mon2,addr_accbuf_mon3,busy,lastshotdone,shotcnt,test1,procdone,cnt00,cnt01,cnt02,cnt03,cnt10,cnt11,cnt12,cnt13,cnt20,cnt21,cnt22,cnt23,cnt30,cnt31,cnt32,cnt33,addr_sdbuf_mon0,addr_sdbuf_mon1
);
logic [DATA_WIDTH-1:0] rdata;
logic [DATA_WIDTH-1:0] wdata;
logic [ADDR_WIDTH-1:0] waddr;
logic [1-1:0] wren;

wire [32-1:0] resetacc;reg [32-1:0] reg_resetacc=0;reg stb_resetacc;assign resetacc=reg_resetacc;
wire [32-1:0] addr_accbuf_mon0;
wire [32-1:0] addr_accbuf_mon1;
wire [32-1:0] addr_accbuf_mon2;
wire [32-1:0] addr_accbuf_mon3;
wire [32-1:0] amp;reg [32-1:0] reg_amp=32000;reg stb_amp;assign amp=reg_amp;
wire [32-1:0] bramsel;reg [32-1:0] reg_bramsel=0;reg stb_bramsel;assign bramsel=reg_bramsel;
wire [4-1:0] busy;
wire [32-1:0] coef00;reg [32-1:0] reg_coef00=2147418112;reg stb_coef00;assign coef00=reg_coef00;
wire [32-1:0] coef01;reg [32-1:0] reg_coef01=0;reg stb_coef01;assign coef01=reg_coef01;
wire [32-1:0] coef02;reg [32-1:0] reg_coef02=0;reg stb_coef02;assign coef02=reg_coef02;
wire [32-1:0] coef03;reg [32-1:0] reg_coef03=0;reg stb_coef03;assign coef03=reg_coef03;
wire [32-1:0] coef10;reg [32-1:0] reg_coef10=0;reg stb_coef10;assign coef10=reg_coef10;
wire [32-1:0] coef11;reg [32-1:0] reg_coef11=2147418112;reg stb_coef11;assign coef11=reg_coef11;
wire [32-1:0] coef12;reg [32-1:0] reg_coef12=0;reg stb_coef12;assign coef12=reg_coef12;
wire [32-1:0] coef13;reg [32-1:0] reg_coef13=0;reg stb_coef13;assign coef13=reg_coef13;
wire [32-1:0] coef20;reg [32-1:0] reg_coef20=0;reg stb_coef20;assign coef20=reg_coef20;
wire [32-1:0] coef21;reg [32-1:0] reg_coef21=0;reg stb_coef21;assign coef21=reg_coef21;
wire [32-1:0] coef22;reg [32-1:0] reg_coef22=2147418112;reg stb_coef22;assign coef22=reg_coef22;
wire [32-1:0] coef23;reg [32-1:0] reg_coef23=0;reg stb_coef23;assign coef23=reg_coef23;
wire [32-1:0] coef30;reg [32-1:0] reg_coef30=0;reg stb_coef30;assign coef30=reg_coef30;
wire [32-1:0] coef31;reg [32-1:0] reg_coef31=0;reg stb_coef31;assign coef31=reg_coef31;
wire [32-1:0] coef32;reg [32-1:0] reg_coef32=0;reg stb_coef32;assign coef32=reg_coef32;
wire [32-1:0] coef33;reg [32-1:0] reg_coef33=2147418112;reg stb_coef33;assign coef33=reg_coef33;
wire [32-1:0] dacsel;reg [32-1:0] reg_dacsel=3;reg stb_dacsel;assign dacsel=reg_dacsel;
wire [1-1:0] dspreset;reg [1-1:0] reg_dspreset=0;reg stb_dspreset;assign dspreset=reg_dspreset;
wire [1-1:0] lastshotdone;
wire [32-1:0] nshot;reg [32-1:0] reg_nshot=10;reg stb_nshot;assign nshot=reg_nshot;
wire [32-1:0] qdrvfreqsel;reg [32-1:0] reg_qdrvfreqsel=3;reg stb_qdrvfreqsel;assign qdrvfreqsel=reg_qdrvfreqsel;
wire [32-1:0] rdlofreqsel;reg [32-1:0] reg_rdlofreqsel=3;reg stb_rdlofreqsel;assign rdlofreqsel=reg_rdlofreqsel;
wire [32-1:0] rdrvfreqsel;reg [32-1:0] reg_rdrvfreqsel=3;reg stb_rdrvfreqsel;assign rdrvfreqsel=reg_rdrvfreqsel;
wire [32-1:0] reset_bram_read;reg [32-1:0] reg_reset_bram_read=0;reg stb_reset_bram_read;assign reset_bram_read=reg_reset_bram_read;
wire [32-1:0] shotcnt;
wire [1-1:0] start;reg [1-1:0] reg_start=0;reg stb_start;assign start=reg_start;
wire [32-1:0] test;reg [32-1:0] reg_test=0;reg stb_test;assign test=reg_test;
wire [32-1:0] test1;
wire [1-1:0] acqbufreset;reg [1-1:0] reg_acqbufreset=1;reg stb_acqbufreset;assign acqbufreset=reg_acqbufreset;
wire [1-1:0] dacmonreset;reg [1-1:0] reg_dacmonreset=1;reg stb_dacmonreset;assign dacmonreset=reg_dacmonreset;
wire [8-1:0] decimator;reg [8-1:0] reg_decimator=1;reg stb_decimator;assign decimator=reg_decimator;
wire [5-1:0] acqchansel0;reg [5-1:0] reg_acqchansel0=1;reg stb_acqchansel0;assign acqchansel0=reg_acqchansel0;
wire [5-1:0] acqchansel1;reg [5-1:0] reg_acqchansel1=0;reg stb_acqchansel1;assign acqchansel1=reg_acqchansel1;
wire [5-1:0] dacmonchansel0;reg [5-1:0] reg_dacmonchansel0=0;reg stb_dacmonchansel0;assign dacmonchansel0=reg_dacmonchansel0;
wire [5-1:0] dacmonchansel1;reg [5-1:0] reg_dacmonchansel1=0;reg stb_dacmonchansel1;assign dacmonchansel1=reg_dacmonchansel1;
wire [5-1:0] dacmonchansel2;reg [5-1:0] reg_dacmonchansel2=0;reg stb_dacmonchansel2;assign dacmonchansel2=reg_dacmonchansel2;
wire [5-1:0] dacmonchansel3;reg [5-1:0] reg_dacmonchansel3=0;reg stb_dacmonchansel3;assign dacmonchansel3=reg_dacmonchansel3;
wire [16-1:0] delayaftertrig;reg [16-1:0] reg_delayaftertrig=100;reg stb_delayaftertrig;assign delayaftertrig=reg_delayaftertrig;
wire [16-1:0] mixbb1sel;reg [16-1:0] reg_mixbb1sel=0;reg stb_mixbb1sel;assign mixbb1sel=reg_mixbb1sel;
wire [16-1:0] mixbb2sel;reg [16-1:0] reg_mixbb2sel=1;reg stb_mixbb2sel;assign mixbb2sel=reg_mixbb2sel;
wire [5-1:0] shift;reg [5-1:0] reg_shift=15;reg stb_shift;assign shift=reg_shift;
wire [32-1:0] procdone;
wire [32-1:0] cnt00;
wire [32-1:0] cnt01;
wire [32-1:0] cnt02;
wire [32-1:0] cnt03;
wire [32-1:0] cnt10;
wire [32-1:0] cnt11;
wire [32-1:0] cnt12;
wire [32-1:0] cnt13;
wire [32-1:0] cnt20;
wire [32-1:0] cnt21;
wire [32-1:0] cnt22;
wire [32-1:0] cnt23;
wire [32-1:0] cnt30;
wire [32-1:0] cnt31;
wire [32-1:0] cnt32;
wire [32-1:0] cnt33;
wire [32-1:0] addr_sdbuf_mon0;
wire [32-1:0] addr_sdbuf_mon1;
wire signed [18-1:0] W_Q0_0_0_0;reg signed [18-1:0] reg_W_Q0_0_0_0=65248;reg stb_W_Q0_0_0_0;assign W_Q0_0_0_0=reg_W_Q0_0_0_0;
wire signed [18-1:0] W_Q0_0_0_1;reg signed [18-1:0] reg_W_Q0_0_0_1=65288;reg stb_W_Q0_0_0_1;assign W_Q0_0_0_1=reg_W_Q0_0_0_1;
wire signed [18-1:0] W_Q0_0_0_2;reg signed [18-1:0] reg_W_Q0_0_0_2=65031;reg stb_W_Q0_0_0_2;assign W_Q0_0_0_2=reg_W_Q0_0_0_2;
wire signed [18-1:0] W_Q0_0_0_3;reg signed [18-1:0] reg_W_Q0_0_0_3=346;reg stb_W_Q0_0_0_3;assign W_Q0_0_0_3=reg_W_Q0_0_0_3;
wire signed [18-1:0] W_Q0_0_0_4;reg signed [18-1:0] reg_W_Q0_0_0_4=405;reg stb_W_Q0_0_0_4;assign W_Q0_0_0_4=reg_W_Q0_0_0_4;
wire signed [18-1:0] W_Q0_0_0_5;reg signed [18-1:0] reg_W_Q0_0_0_5=509;reg stb_W_Q0_0_0_5;assign W_Q0_0_0_5=reg_W_Q0_0_0_5;
wire signed [18-1:0] W_Q0_0_0_6;reg signed [18-1:0] reg_W_Q0_0_0_6=869;reg stb_W_Q0_0_0_6;assign W_Q0_0_0_6=reg_W_Q0_0_0_6;
wire signed [18-1:0] W_Q0_0_0_7;reg signed [18-1:0] reg_W_Q0_0_0_7=581;reg stb_W_Q0_0_0_7;assign W_Q0_0_0_7=reg_W_Q0_0_0_7;
wire signed [18-1:0] W_Q0_0_1_0;reg signed [18-1:0] reg_W_Q0_0_1_0=304;reg stb_W_Q0_0_1_0;assign W_Q0_0_1_0=reg_W_Q0_0_1_0;
wire signed [18-1:0] W_Q0_0_1_1;reg signed [18-1:0] reg_W_Q0_0_1_1=65043;reg stb_W_Q0_0_1_1;assign W_Q0_0_1_1=reg_W_Q0_0_1_1;
wire signed [18-1:0] W_Q0_0_1_2;reg signed [18-1:0] reg_W_Q0_0_1_2=65242;reg stb_W_Q0_0_1_2;assign W_Q0_0_1_2=reg_W_Q0_0_1_2;
wire signed [18-1:0] W_Q0_0_1_3;reg signed [18-1:0] reg_W_Q0_0_1_3=319;reg stb_W_Q0_0_1_3;assign W_Q0_0_1_3=reg_W_Q0_0_1_3;
wire signed [18-1:0] W_Q0_0_1_4;reg signed [18-1:0] reg_W_Q0_0_1_4=64877;reg stb_W_Q0_0_1_4;assign W_Q0_0_1_4=reg_W_Q0_0_1_4;
wire signed [18-1:0] W_Q0_0_1_5;reg signed [18-1:0] reg_W_Q0_0_1_5=124;reg stb_W_Q0_0_1_5;assign W_Q0_0_1_5=reg_W_Q0_0_1_5;
wire signed [18-1:0] W_Q0_0_1_6;reg signed [18-1:0] reg_W_Q0_0_1_6=65192;reg stb_W_Q0_0_1_6;assign W_Q0_0_1_6=reg_W_Q0_0_1_6;
wire signed [18-1:0] W_Q0_0_1_7;reg signed [18-1:0] reg_W_Q0_0_1_7=65348;reg stb_W_Q0_0_1_7;assign W_Q0_0_1_7=reg_W_Q0_0_1_7;
wire signed [18-1:0] W_Q0_1_0_0;reg signed [18-1:0] reg_W_Q0_1_0_0=394;reg stb_W_Q0_1_0_0;assign W_Q0_1_0_0=reg_W_Q0_1_0_0;
wire signed [18-1:0] W_Q0_1_0_1;reg signed [18-1:0] reg_W_Q0_1_0_1=65201;reg stb_W_Q0_1_0_1;assign W_Q0_1_0_1=reg_W_Q0_1_0_1;
wire signed [18-1:0] W_Q0_1_0_2;reg signed [18-1:0] reg_W_Q0_1_0_2=943;reg stb_W_Q0_1_0_2;assign W_Q0_1_0_2=reg_W_Q0_1_0_2;
wire signed [18-1:0] W_Q0_1_0_3;reg signed [18-1:0] reg_W_Q0_1_0_3=65470;reg stb_W_Q0_1_0_3;assign W_Q0_1_0_3=reg_W_Q0_1_0_3;
wire signed [18-1:0] W_Q0_1_1_0;reg signed [18-1:0] reg_W_Q0_1_1_0=642;reg stb_W_Q0_1_1_0;assign W_Q0_1_1_0=reg_W_Q0_1_1_0;
wire signed [18-1:0] W_Q0_1_1_1;reg signed [18-1:0] reg_W_Q0_1_1_1=44;reg stb_W_Q0_1_1_1;assign W_Q0_1_1_1=reg_W_Q0_1_1_1;
wire signed [18-1:0] W_Q0_1_1_2;reg signed [18-1:0] reg_W_Q0_1_1_2=64664;reg stb_W_Q0_1_1_2;assign W_Q0_1_1_2=reg_W_Q0_1_1_2;
wire signed [18-1:0] W_Q0_1_1_3;reg signed [18-1:0] reg_W_Q0_1_1_3=718;reg stb_W_Q0_1_1_3;assign W_Q0_1_1_3=reg_W_Q0_1_1_3;
wire signed [18-1:0] W_Q0_1_2_0;reg signed [18-1:0] reg_W_Q0_1_2_0=172;reg stb_W_Q0_1_2_0;assign W_Q0_1_2_0=reg_W_Q0_1_2_0;
wire signed [18-1:0] W_Q0_1_2_1;reg signed [18-1:0] reg_W_Q0_1_2_1=65162;reg stb_W_Q0_1_2_1;assign W_Q0_1_2_1=reg_W_Q0_1_2_1;
wire signed [18-1:0] W_Q0_1_2_2;reg signed [18-1:0] reg_W_Q0_1_2_2=700;reg stb_W_Q0_1_2_2;assign W_Q0_1_2_2=reg_W_Q0_1_2_2;
wire signed [18-1:0] W_Q0_1_2_3;reg signed [18-1:0] reg_W_Q0_1_2_3=828;reg stb_W_Q0_1_2_3;assign W_Q0_1_2_3=reg_W_Q0_1_2_3;
wire signed [18-1:0] W_Q0_1_3_0;reg signed [18-1:0] reg_W_Q0_1_3_0=202;reg stb_W_Q0_1_3_0;assign W_Q0_1_3_0=reg_W_Q0_1_3_0;
wire signed [18-1:0] W_Q0_1_3_1;reg signed [18-1:0] reg_W_Q0_1_3_1=65060;reg stb_W_Q0_1_3_1;assign W_Q0_1_3_1=reg_W_Q0_1_3_1;
wire signed [18-1:0] W_Q0_1_3_2;reg signed [18-1:0] reg_W_Q0_1_3_2=1179;reg stb_W_Q0_1_3_2;assign W_Q0_1_3_2=reg_W_Q0_1_3_2;
wire signed [18-1:0] W_Q0_1_3_3;reg signed [18-1:0] reg_W_Q0_1_3_3=64947;reg stb_W_Q0_1_3_3;assign W_Q0_1_3_3=reg_W_Q0_1_3_3;
wire signed [18-1:0] W_Q0_1_4_0;reg signed [18-1:0] reg_W_Q0_1_4_0=10;reg stb_W_Q0_1_4_0;assign W_Q0_1_4_0=reg_W_Q0_1_4_0;
wire signed [18-1:0] W_Q0_1_4_1;reg signed [18-1:0] reg_W_Q0_1_4_1=704;reg stb_W_Q0_1_4_1;assign W_Q0_1_4_1=reg_W_Q0_1_4_1;
wire signed [18-1:0] W_Q0_1_4_2;reg signed [18-1:0] reg_W_Q0_1_4_2=65402;reg stb_W_Q0_1_4_2;assign W_Q0_1_4_2=reg_W_Q0_1_4_2;
wire signed [18-1:0] W_Q0_1_4_3;reg signed [18-1:0] reg_W_Q0_1_4_3=65316;reg stb_W_Q0_1_4_3;assign W_Q0_1_4_3=reg_W_Q0_1_4_3;
wire signed [18-1:0] W_Q0_1_5_0;reg signed [18-1:0] reg_W_Q0_1_5_0=330;reg stb_W_Q0_1_5_0;assign W_Q0_1_5_0=reg_W_Q0_1_5_0;
wire signed [18-1:0] W_Q0_1_5_1;reg signed [18-1:0] reg_W_Q0_1_5_1=64795;reg stb_W_Q0_1_5_1;assign W_Q0_1_5_1=reg_W_Q0_1_5_1;
wire signed [18-1:0] W_Q0_1_5_2;reg signed [18-1:0] reg_W_Q0_1_5_2=432;reg stb_W_Q0_1_5_2;assign W_Q0_1_5_2=reg_W_Q0_1_5_2;
wire signed [18-1:0] W_Q0_1_5_3;reg signed [18-1:0] reg_W_Q0_1_5_3=37;reg stb_W_Q0_1_5_3;assign W_Q0_1_5_3=reg_W_Q0_1_5_3;
wire signed [18-1:0] W_Q0_1_6_0;reg signed [18-1:0] reg_W_Q0_1_6_0=64817;reg stb_W_Q0_1_6_0;assign W_Q0_1_6_0=reg_W_Q0_1_6_0;
wire signed [18-1:0] W_Q0_1_6_1;reg signed [18-1:0] reg_W_Q0_1_6_1=65506;reg stb_W_Q0_1_6_1;assign W_Q0_1_6_1=reg_W_Q0_1_6_1;
wire signed [18-1:0] W_Q0_1_6_2;reg signed [18-1:0] reg_W_Q0_1_6_2=70;reg stb_W_Q0_1_6_2;assign W_Q0_1_6_2=reg_W_Q0_1_6_2;
wire signed [18-1:0] W_Q0_1_6_3;reg signed [18-1:0] reg_W_Q0_1_6_3=65507;reg stb_W_Q0_1_6_3;assign W_Q0_1_6_3=reg_W_Q0_1_6_3;
wire signed [18-1:0] W_Q0_1_7_0;reg signed [18-1:0] reg_W_Q0_1_7_0=302;reg stb_W_Q0_1_7_0;assign W_Q0_1_7_0=reg_W_Q0_1_7_0;
wire signed [18-1:0] W_Q0_1_7_1;reg signed [18-1:0] reg_W_Q0_1_7_1=65497;reg stb_W_Q0_1_7_1;assign W_Q0_1_7_1=reg_W_Q0_1_7_1;
wire signed [18-1:0] W_Q0_1_7_2;reg signed [18-1:0] reg_W_Q0_1_7_2=200;reg stb_W_Q0_1_7_2;assign W_Q0_1_7_2=reg_W_Q0_1_7_2;
wire signed [18-1:0] W_Q0_1_7_3;reg signed [18-1:0] reg_W_Q0_1_7_3=145;reg stb_W_Q0_1_7_3;assign W_Q0_1_7_3=reg_W_Q0_1_7_3;
wire signed [18-1:0] W_Q0_2_0_0;reg signed [18-1:0] reg_W_Q0_2_0_0=64822;reg stb_W_Q0_2_0_0;assign W_Q0_2_0_0=reg_W_Q0_2_0_0;
wire signed [18-1:0] W_Q0_2_1_0;reg signed [18-1:0] reg_W_Q0_2_1_0=65139;reg stb_W_Q0_2_1_0;assign W_Q0_2_1_0=reg_W_Q0_2_1_0;
wire signed [18-1:0] W_Q0_2_2_0;reg signed [18-1:0] reg_W_Q0_2_2_0=911;reg stb_W_Q0_2_2_0;assign W_Q0_2_2_0=reg_W_Q0_2_2_0;
wire signed [18-1:0] W_Q0_2_3_0;reg signed [18-1:0] reg_W_Q0_2_3_0=64698;reg stb_W_Q0_2_3_0;assign W_Q0_2_3_0=reg_W_Q0_2_3_0;
wire signed [18-1:0] B_Q0_0_0;reg signed [18-1:0] reg_B_Q0_0_0=157;reg stb_B_Q0_0_0;assign B_Q0_0_0=reg_B_Q0_0_0;
wire signed [18-1:0] B_Q0_0_1;reg signed [18-1:0] reg_B_Q0_0_1=111;reg stb_B_Q0_0_1;assign B_Q0_0_1=reg_B_Q0_0_1;
wire signed [18-1:0] B_Q0_0_2;reg signed [18-1:0] reg_B_Q0_0_2=240;reg stb_B_Q0_0_2;assign B_Q0_0_2=reg_B_Q0_0_2;
wire signed [18-1:0] B_Q0_0_3;reg signed [18-1:0] reg_B_Q0_0_3=325;reg stb_B_Q0_0_3;assign B_Q0_0_3=reg_B_Q0_0_3;
wire signed [18-1:0] B_Q0_0_4;reg signed [18-1:0] reg_B_Q0_0_4=65370;reg stb_B_Q0_0_4;assign B_Q0_0_4=reg_B_Q0_0_4;
wire signed [18-1:0] B_Q0_0_5;reg signed [18-1:0] reg_B_Q0_0_5=65487;reg stb_B_Q0_0_5;assign B_Q0_0_5=reg_B_Q0_0_5;
wire signed [18-1:0] B_Q0_0_6;reg signed [18-1:0] reg_B_Q0_0_6=38;reg stb_B_Q0_0_6;assign B_Q0_0_6=reg_B_Q0_0_6;
wire signed [18-1:0] B_Q0_0_7;reg signed [18-1:0] reg_B_Q0_0_7=65448;reg stb_B_Q0_0_7;assign B_Q0_0_7=reg_B_Q0_0_7;
wire signed [18-1:0] B_Q0_1_0;reg signed [18-1:0] reg_B_Q0_1_0=65260;reg stb_B_Q0_1_0;assign B_Q0_1_0=reg_B_Q0_1_0;
wire signed [18-1:0] B_Q0_1_1;reg signed [18-1:0] reg_B_Q0_1_1=159;reg stb_B_Q0_1_1;assign B_Q0_1_1=reg_B_Q0_1_1;
wire signed [18-1:0] B_Q0_1_2;reg signed [18-1:0] reg_B_Q0_1_2=358;reg stb_B_Q0_1_2;assign B_Q0_1_2=reg_B_Q0_1_2;
wire signed [18-1:0] B_Q0_1_3;reg signed [18-1:0] reg_B_Q0_1_3=65423;reg stb_B_Q0_1_3;assign B_Q0_1_3=reg_B_Q0_1_3;
wire signed [18-1:0] B_Q0_2_0;reg signed [18-1:0] reg_B_Q0_2_0=333;reg stb_B_Q0_2_0;assign B_Q0_2_0=reg_B_Q0_2_0;
wire signed [18-1:0] W_Q1_0_0_0;reg signed [18-1:0] reg_W_Q1_0_0_0=65248;reg stb_W_Q1_0_0_0;assign W_Q1_0_0_0=reg_W_Q1_0_0_0;
wire signed [18-1:0] W_Q1_0_0_1;reg signed [18-1:0] reg_W_Q1_0_0_1=65288;reg stb_W_Q1_0_0_1;assign W_Q1_0_0_1=reg_W_Q1_0_0_1;
wire signed [18-1:0] W_Q1_0_0_2;reg signed [18-1:0] reg_W_Q1_0_0_2=65031;reg stb_W_Q1_0_0_2;assign W_Q1_0_0_2=reg_W_Q1_0_0_2;
wire signed [18-1:0] W_Q1_0_0_3;reg signed [18-1:0] reg_W_Q1_0_0_3=346;reg stb_W_Q1_0_0_3;assign W_Q1_0_0_3=reg_W_Q1_0_0_3;
wire signed [18-1:0] W_Q1_0_0_4;reg signed [18-1:0] reg_W_Q1_0_0_4=405;reg stb_W_Q1_0_0_4;assign W_Q1_0_0_4=reg_W_Q1_0_0_4;
wire signed [18-1:0] W_Q1_0_0_5;reg signed [18-1:0] reg_W_Q1_0_0_5=509;reg stb_W_Q1_0_0_5;assign W_Q1_0_0_5=reg_W_Q1_0_0_5;
wire signed [18-1:0] W_Q1_0_0_6;reg signed [18-1:0] reg_W_Q1_0_0_6=869;reg stb_W_Q1_0_0_6;assign W_Q1_0_0_6=reg_W_Q1_0_0_6;
wire signed [18-1:0] W_Q1_0_0_7;reg signed [18-1:0] reg_W_Q1_0_0_7=581;reg stb_W_Q1_0_0_7;assign W_Q1_0_0_7=reg_W_Q1_0_0_7;
wire signed [18-1:0] W_Q1_0_1_0;reg signed [18-1:0] reg_W_Q1_0_1_0=304;reg stb_W_Q1_0_1_0;assign W_Q1_0_1_0=reg_W_Q1_0_1_0;
wire signed [18-1:0] W_Q1_0_1_1;reg signed [18-1:0] reg_W_Q1_0_1_1=65043;reg stb_W_Q1_0_1_1;assign W_Q1_0_1_1=reg_W_Q1_0_1_1;
wire signed [18-1:0] W_Q1_0_1_2;reg signed [18-1:0] reg_W_Q1_0_1_2=65242;reg stb_W_Q1_0_1_2;assign W_Q1_0_1_2=reg_W_Q1_0_1_2;
wire signed [18-1:0] W_Q1_0_1_3;reg signed [18-1:0] reg_W_Q1_0_1_3=319;reg stb_W_Q1_0_1_3;assign W_Q1_0_1_3=reg_W_Q1_0_1_3;
wire signed [18-1:0] W_Q1_0_1_4;reg signed [18-1:0] reg_W_Q1_0_1_4=64877;reg stb_W_Q1_0_1_4;assign W_Q1_0_1_4=reg_W_Q1_0_1_4;
wire signed [18-1:0] W_Q1_0_1_5;reg signed [18-1:0] reg_W_Q1_0_1_5=124;reg stb_W_Q1_0_1_5;assign W_Q1_0_1_5=reg_W_Q1_0_1_5;
wire signed [18-1:0] W_Q1_0_1_6;reg signed [18-1:0] reg_W_Q1_0_1_6=65192;reg stb_W_Q1_0_1_6;assign W_Q1_0_1_6=reg_W_Q1_0_1_6;
wire signed [18-1:0] W_Q1_0_1_7;reg signed [18-1:0] reg_W_Q1_0_1_7=65348;reg stb_W_Q1_0_1_7;assign W_Q1_0_1_7=reg_W_Q1_0_1_7;
wire signed [18-1:0] W_Q1_1_0_0;reg signed [18-1:0] reg_W_Q1_1_0_0=394;reg stb_W_Q1_1_0_0;assign W_Q1_1_0_0=reg_W_Q1_1_0_0;
wire signed [18-1:0] W_Q1_1_0_1;reg signed [18-1:0] reg_W_Q1_1_0_1=65201;reg stb_W_Q1_1_0_1;assign W_Q1_1_0_1=reg_W_Q1_1_0_1;
wire signed [18-1:0] W_Q1_1_0_2;reg signed [18-1:0] reg_W_Q1_1_0_2=943;reg stb_W_Q1_1_0_2;assign W_Q1_1_0_2=reg_W_Q1_1_0_2;
wire signed [18-1:0] W_Q1_1_0_3;reg signed [18-1:0] reg_W_Q1_1_0_3=65470;reg stb_W_Q1_1_0_3;assign W_Q1_1_0_3=reg_W_Q1_1_0_3;
wire signed [18-1:0] W_Q1_1_1_0;reg signed [18-1:0] reg_W_Q1_1_1_0=642;reg stb_W_Q1_1_1_0;assign W_Q1_1_1_0=reg_W_Q1_1_1_0;
wire signed [18-1:0] W_Q1_1_1_1;reg signed [18-1:0] reg_W_Q1_1_1_1=44;reg stb_W_Q1_1_1_1;assign W_Q1_1_1_1=reg_W_Q1_1_1_1;
wire signed [18-1:0] W_Q1_1_1_2;reg signed [18-1:0] reg_W_Q1_1_1_2=64664;reg stb_W_Q1_1_1_2;assign W_Q1_1_1_2=reg_W_Q1_1_1_2;
wire signed [18-1:0] W_Q1_1_1_3;reg signed [18-1:0] reg_W_Q1_1_1_3=718;reg stb_W_Q1_1_1_3;assign W_Q1_1_1_3=reg_W_Q1_1_1_3;
wire signed [18-1:0] W_Q1_1_2_0;reg signed [18-1:0] reg_W_Q1_1_2_0=172;reg stb_W_Q1_1_2_0;assign W_Q1_1_2_0=reg_W_Q1_1_2_0;
wire signed [18-1:0] W_Q1_1_2_1;reg signed [18-1:0] reg_W_Q1_1_2_1=65162;reg stb_W_Q1_1_2_1;assign W_Q1_1_2_1=reg_W_Q1_1_2_1;
wire signed [18-1:0] W_Q1_1_2_2;reg signed [18-1:0] reg_W_Q1_1_2_2=700;reg stb_W_Q1_1_2_2;assign W_Q1_1_2_2=reg_W_Q1_1_2_2;
wire signed [18-1:0] W_Q1_1_2_3;reg signed [18-1:0] reg_W_Q1_1_2_3=828;reg stb_W_Q1_1_2_3;assign W_Q1_1_2_3=reg_W_Q1_1_2_3;
wire signed [18-1:0] W_Q1_1_3_0;reg signed [18-1:0] reg_W_Q1_1_3_0=202;reg stb_W_Q1_1_3_0;assign W_Q1_1_3_0=reg_W_Q1_1_3_0;
wire signed [18-1:0] W_Q1_1_3_1;reg signed [18-1:0] reg_W_Q1_1_3_1=65060;reg stb_W_Q1_1_3_1;assign W_Q1_1_3_1=reg_W_Q1_1_3_1;
wire signed [18-1:0] W_Q1_1_3_2;reg signed [18-1:0] reg_W_Q1_1_3_2=1179;reg stb_W_Q1_1_3_2;assign W_Q1_1_3_2=reg_W_Q1_1_3_2;
wire signed [18-1:0] W_Q1_1_3_3;reg signed [18-1:0] reg_W_Q1_1_3_3=64947;reg stb_W_Q1_1_3_3;assign W_Q1_1_3_3=reg_W_Q1_1_3_3;
wire signed [18-1:0] W_Q1_1_4_0;reg signed [18-1:0] reg_W_Q1_1_4_0=10;reg stb_W_Q1_1_4_0;assign W_Q1_1_4_0=reg_W_Q1_1_4_0;
wire signed [18-1:0] W_Q1_1_4_1;reg signed [18-1:0] reg_W_Q1_1_4_1=704;reg stb_W_Q1_1_4_1;assign W_Q1_1_4_1=reg_W_Q1_1_4_1;
wire signed [18-1:0] W_Q1_1_4_2;reg signed [18-1:0] reg_W_Q1_1_4_2=65402;reg stb_W_Q1_1_4_2;assign W_Q1_1_4_2=reg_W_Q1_1_4_2;
wire signed [18-1:0] W_Q1_1_4_3;reg signed [18-1:0] reg_W_Q1_1_4_3=65316;reg stb_W_Q1_1_4_3;assign W_Q1_1_4_3=reg_W_Q1_1_4_3;
wire signed [18-1:0] W_Q1_1_5_0;reg signed [18-1:0] reg_W_Q1_1_5_0=330;reg stb_W_Q1_1_5_0;assign W_Q1_1_5_0=reg_W_Q1_1_5_0;
wire signed [18-1:0] W_Q1_1_5_1;reg signed [18-1:0] reg_W_Q1_1_5_1=64795;reg stb_W_Q1_1_5_1;assign W_Q1_1_5_1=reg_W_Q1_1_5_1;
wire signed [18-1:0] W_Q1_1_5_2;reg signed [18-1:0] reg_W_Q1_1_5_2=432;reg stb_W_Q1_1_5_2;assign W_Q1_1_5_2=reg_W_Q1_1_5_2;
wire signed [18-1:0] W_Q1_1_5_3;reg signed [18-1:0] reg_W_Q1_1_5_3=37;reg stb_W_Q1_1_5_3;assign W_Q1_1_5_3=reg_W_Q1_1_5_3;
wire signed [18-1:0] W_Q1_1_6_0;reg signed [18-1:0] reg_W_Q1_1_6_0=64817;reg stb_W_Q1_1_6_0;assign W_Q1_1_6_0=reg_W_Q1_1_6_0;
wire signed [18-1:0] W_Q1_1_6_1;reg signed [18-1:0] reg_W_Q1_1_6_1=65506;reg stb_W_Q1_1_6_1;assign W_Q1_1_6_1=reg_W_Q1_1_6_1;
wire signed [18-1:0] W_Q1_1_6_2;reg signed [18-1:0] reg_W_Q1_1_6_2=70;reg stb_W_Q1_1_6_2;assign W_Q1_1_6_2=reg_W_Q1_1_6_2;
wire signed [18-1:0] W_Q1_1_6_3;reg signed [18-1:0] reg_W_Q1_1_6_3=65507;reg stb_W_Q1_1_6_3;assign W_Q1_1_6_3=reg_W_Q1_1_6_3;
wire signed [18-1:0] W_Q1_1_7_0;reg signed [18-1:0] reg_W_Q1_1_7_0=302;reg stb_W_Q1_1_7_0;assign W_Q1_1_7_0=reg_W_Q1_1_7_0;
wire signed [18-1:0] W_Q1_1_7_1;reg signed [18-1:0] reg_W_Q1_1_7_1=65497;reg stb_W_Q1_1_7_1;assign W_Q1_1_7_1=reg_W_Q1_1_7_1;
wire signed [18-1:0] W_Q1_1_7_2;reg signed [18-1:0] reg_W_Q1_1_7_2=200;reg stb_W_Q1_1_7_2;assign W_Q1_1_7_2=reg_W_Q1_1_7_2;
wire signed [18-1:0] W_Q1_1_7_3;reg signed [18-1:0] reg_W_Q1_1_7_3=145;reg stb_W_Q1_1_7_3;assign W_Q1_1_7_3=reg_W_Q1_1_7_3;
wire signed [18-1:0] W_Q1_2_0_0;reg signed [18-1:0] reg_W_Q1_2_0_0=64822;reg stb_W_Q1_2_0_0;assign W_Q1_2_0_0=reg_W_Q1_2_0_0;
wire signed [18-1:0] W_Q1_2_1_0;reg signed [18-1:0] reg_W_Q1_2_1_0=65139;reg stb_W_Q1_2_1_0;assign W_Q1_2_1_0=reg_W_Q1_2_1_0;
wire signed [18-1:0] W_Q1_2_2_0;reg signed [18-1:0] reg_W_Q1_2_2_0=911;reg stb_W_Q1_2_2_0;assign W_Q1_2_2_0=reg_W_Q1_2_2_0;
wire signed [18-1:0] W_Q1_2_3_0;reg signed [18-1:0] reg_W_Q1_2_3_0=64698;reg stb_W_Q1_2_3_0;assign W_Q1_2_3_0=reg_W_Q1_2_3_0;
wire signed [18-1:0] B_Q1_0_0;reg signed [18-1:0] reg_B_Q1_0_0=157;reg stb_B_Q1_0_0;assign B_Q1_0_0=reg_B_Q1_0_0;
wire signed [18-1:0] B_Q1_0_1;reg signed [18-1:0] reg_B_Q1_0_1=111;reg stb_B_Q1_0_1;assign B_Q1_0_1=reg_B_Q1_0_1;
wire signed [18-1:0] B_Q1_0_2;reg signed [18-1:0] reg_B_Q1_0_2=240;reg stb_B_Q1_0_2;assign B_Q1_0_2=reg_B_Q1_0_2;
wire signed [18-1:0] B_Q1_0_3;reg signed [18-1:0] reg_B_Q1_0_3=325;reg stb_B_Q1_0_3;assign B_Q1_0_3=reg_B_Q1_0_3;
wire signed [18-1:0] B_Q1_0_4;reg signed [18-1:0] reg_B_Q1_0_4=65370;reg stb_B_Q1_0_4;assign B_Q1_0_4=reg_B_Q1_0_4;
wire signed [18-1:0] B_Q1_0_5;reg signed [18-1:0] reg_B_Q1_0_5=65487;reg stb_B_Q1_0_5;assign B_Q1_0_5=reg_B_Q1_0_5;
wire signed [18-1:0] B_Q1_0_6;reg signed [18-1:0] reg_B_Q1_0_6=38;reg stb_B_Q1_0_6;assign B_Q1_0_6=reg_B_Q1_0_6;
wire signed [18-1:0] B_Q1_0_7;reg signed [18-1:0] reg_B_Q1_0_7=65448;reg stb_B_Q1_0_7;assign B_Q1_0_7=reg_B_Q1_0_7;
wire signed [18-1:0] B_Q1_1_0;reg signed [18-1:0] reg_B_Q1_1_0=65260;reg stb_B_Q1_1_0;assign B_Q1_1_0=reg_B_Q1_1_0;
wire signed [18-1:0] B_Q1_1_1;reg signed [18-1:0] reg_B_Q1_1_1=159;reg stb_B_Q1_1_1;assign B_Q1_1_1=reg_B_Q1_1_1;
wire signed [18-1:0] B_Q1_1_2;reg signed [18-1:0] reg_B_Q1_1_2=358;reg stb_B_Q1_1_2;assign B_Q1_1_2=reg_B_Q1_1_2;
wire signed [18-1:0] B_Q1_1_3;reg signed [18-1:0] reg_B_Q1_1_3=65423;reg stb_B_Q1_1_3;assign B_Q1_1_3=reg_B_Q1_1_3;
wire signed [18-1:0] B_Q1_2_0;reg signed [18-1:0] reg_B_Q1_2_0=333;reg stb_B_Q1_2_0;assign B_Q1_2_0=reg_B_Q1_2_0;
wire signed [18-1:0] W_Q2_0_0_0;reg signed [18-1:0] reg_W_Q2_0_0_0=260183;reg stb_W_Q2_0_0_0;assign W_Q2_0_0_0=reg_W_Q2_0_0_0;
wire signed [18-1:0] W_Q2_0_0_1;reg signed [18-1:0] reg_W_Q2_0_0_1=4862;reg stb_W_Q2_0_0_1;assign W_Q2_0_0_1=reg_W_Q2_0_0_1;
wire signed [18-1:0] W_Q2_0_0_2;reg signed [18-1:0] reg_W_Q2_0_0_2=261334;reg stb_W_Q2_0_0_2;assign W_Q2_0_0_2=reg_W_Q2_0_0_2;
wire signed [18-1:0] W_Q2_0_0_3;reg signed [18-1:0] reg_W_Q2_0_0_3=260711;reg stb_W_Q2_0_0_3;assign W_Q2_0_0_3=reg_W_Q2_0_0_3;
wire signed [18-1:0] W_Q2_0_0_4;reg signed [18-1:0] reg_W_Q2_0_0_4=262141;reg stb_W_Q2_0_0_4;assign W_Q2_0_0_4=reg_W_Q2_0_0_4;
wire signed [18-1:0] W_Q2_0_0_5;reg signed [18-1:0] reg_W_Q2_0_0_5=259938;reg stb_W_Q2_0_0_5;assign W_Q2_0_0_5=reg_W_Q2_0_0_5;
wire signed [18-1:0] W_Q2_0_0_6;reg signed [18-1:0] reg_W_Q2_0_0_6=4215;reg stb_W_Q2_0_0_6;assign W_Q2_0_0_6=reg_W_Q2_0_0_6;
wire signed [18-1:0] W_Q2_0_0_7;reg signed [18-1:0] reg_W_Q2_0_0_7=4895;reg stb_W_Q2_0_0_7;assign W_Q2_0_0_7=reg_W_Q2_0_0_7;
wire signed [18-1:0] W_Q2_0_1_0;reg signed [18-1:0] reg_W_Q2_0_1_0=1258;reg stb_W_Q2_0_1_0;assign W_Q2_0_1_0=reg_W_Q2_0_1_0;
wire signed [18-1:0] W_Q2_0_1_1;reg signed [18-1:0] reg_W_Q2_0_1_1=4406;reg stb_W_Q2_0_1_1;assign W_Q2_0_1_1=reg_W_Q2_0_1_1;
wire signed [18-1:0] W_Q2_0_1_2;reg signed [18-1:0] reg_W_Q2_0_1_2=259194;reg stb_W_Q2_0_1_2;assign W_Q2_0_1_2=reg_W_Q2_0_1_2;
wire signed [18-1:0] W_Q2_0_1_3;reg signed [18-1:0] reg_W_Q2_0_1_3=260609;reg stb_W_Q2_0_1_3;assign W_Q2_0_1_3=reg_W_Q2_0_1_3;
wire signed [18-1:0] W_Q2_0_1_4;reg signed [18-1:0] reg_W_Q2_0_1_4=260881;reg stb_W_Q2_0_1_4;assign W_Q2_0_1_4=reg_W_Q2_0_1_4;
wire signed [18-1:0] W_Q2_0_1_5;reg signed [18-1:0] reg_W_Q2_0_1_5=261883;reg stb_W_Q2_0_1_5;assign W_Q2_0_1_5=reg_W_Q2_0_1_5;
wire signed [18-1:0] W_Q2_0_1_6;reg signed [18-1:0] reg_W_Q2_0_1_6=3074;reg stb_W_Q2_0_1_6;assign W_Q2_0_1_6=reg_W_Q2_0_1_6;
wire signed [18-1:0] W_Q2_0_1_7;reg signed [18-1:0] reg_W_Q2_0_1_7=2106;reg stb_W_Q2_0_1_7;assign W_Q2_0_1_7=reg_W_Q2_0_1_7;
wire signed [18-1:0] W_Q2_1_0_0;reg signed [18-1:0] reg_W_Q2_1_0_0=260105;reg stb_W_Q2_1_0_0;assign W_Q2_1_0_0=reg_W_Q2_1_0_0;
wire signed [18-1:0] W_Q2_1_0_1;reg signed [18-1:0] reg_W_Q2_1_0_1=261076;reg stb_W_Q2_1_0_1;assign W_Q2_1_0_1=reg_W_Q2_1_0_1;
wire signed [18-1:0] W_Q2_1_0_2;reg signed [18-1:0] reg_W_Q2_1_0_2=1240;reg stb_W_Q2_1_0_2;assign W_Q2_1_0_2=reg_W_Q2_1_0_2;
wire signed [18-1:0] W_Q2_1_0_3;reg signed [18-1:0] reg_W_Q2_1_0_3=2377;reg stb_W_Q2_1_0_3;assign W_Q2_1_0_3=reg_W_Q2_1_0_3;
wire signed [18-1:0] W_Q2_1_1_0;reg signed [18-1:0] reg_W_Q2_1_1_0=260362;reg stb_W_Q2_1_1_0;assign W_Q2_1_1_0=reg_W_Q2_1_1_0;
wire signed [18-1:0] W_Q2_1_1_1;reg signed [18-1:0] reg_W_Q2_1_1_1=6050;reg stb_W_Q2_1_1_1;assign W_Q2_1_1_1=reg_W_Q2_1_1_1;
wire signed [18-1:0] W_Q2_1_1_2;reg signed [18-1:0] reg_W_Q2_1_1_2=261792;reg stb_W_Q2_1_1_2;assign W_Q2_1_1_2=reg_W_Q2_1_1_2;
wire signed [18-1:0] W_Q2_1_1_3;reg signed [18-1:0] reg_W_Q2_1_1_3=7072;reg stb_W_Q2_1_1_3;assign W_Q2_1_1_3=reg_W_Q2_1_1_3;
wire signed [18-1:0] W_Q2_1_2_0;reg signed [18-1:0] reg_W_Q2_1_2_0=261219;reg stb_W_Q2_1_2_0;assign W_Q2_1_2_0=reg_W_Q2_1_2_0;
wire signed [18-1:0] W_Q2_1_2_1;reg signed [18-1:0] reg_W_Q2_1_2_1=261083;reg stb_W_Q2_1_2_1;assign W_Q2_1_2_1=reg_W_Q2_1_2_1;
wire signed [18-1:0] W_Q2_1_2_2;reg signed [18-1:0] reg_W_Q2_1_2_2=231;reg stb_W_Q2_1_2_2;assign W_Q2_1_2_2=reg_W_Q2_1_2_2;
wire signed [18-1:0] W_Q2_1_2_3;reg signed [18-1:0] reg_W_Q2_1_2_3=2514;reg stb_W_Q2_1_2_3;assign W_Q2_1_2_3=reg_W_Q2_1_2_3;
wire signed [18-1:0] W_Q2_1_3_0;reg signed [18-1:0] reg_W_Q2_1_3_0=1992;reg stb_W_Q2_1_3_0;assign W_Q2_1_3_0=reg_W_Q2_1_3_0;
wire signed [18-1:0] W_Q2_1_3_1;reg signed [18-1:0] reg_W_Q2_1_3_1=2883;reg stb_W_Q2_1_3_1;assign W_Q2_1_3_1=reg_W_Q2_1_3_1;
wire signed [18-1:0] W_Q2_1_3_2;reg signed [18-1:0] reg_W_Q2_1_3_2=260124;reg stb_W_Q2_1_3_2;assign W_Q2_1_3_2=reg_W_Q2_1_3_2;
wire signed [18-1:0] W_Q2_1_3_3;reg signed [18-1:0] reg_W_Q2_1_3_3=260161;reg stb_W_Q2_1_3_3;assign W_Q2_1_3_3=reg_W_Q2_1_3_3;
wire signed [18-1:0] W_Q2_1_4_0;reg signed [18-1:0] reg_W_Q2_1_4_0=260317;reg stb_W_Q2_1_4_0;assign W_Q2_1_4_0=reg_W_Q2_1_4_0;
wire signed [18-1:0] W_Q2_1_4_1;reg signed [18-1:0] reg_W_Q2_1_4_1=259731;reg stb_W_Q2_1_4_1;assign W_Q2_1_4_1=reg_W_Q2_1_4_1;
wire signed [18-1:0] W_Q2_1_4_2;reg signed [18-1:0] reg_W_Q2_1_4_2=261824;reg stb_W_Q2_1_4_2;assign W_Q2_1_4_2=reg_W_Q2_1_4_2;
wire signed [18-1:0] W_Q2_1_4_3;reg signed [18-1:0] reg_W_Q2_1_4_3=261593;reg stb_W_Q2_1_4_3;assign W_Q2_1_4_3=reg_W_Q2_1_4_3;
wire signed [18-1:0] W_Q2_1_5_0;reg signed [18-1:0] reg_W_Q2_1_5_0=2757;reg stb_W_Q2_1_5_0;assign W_Q2_1_5_0=reg_W_Q2_1_5_0;
wire signed [18-1:0] W_Q2_1_5_1;reg signed [18-1:0] reg_W_Q2_1_5_1=261239;reg stb_W_Q2_1_5_1;assign W_Q2_1_5_1=reg_W_Q2_1_5_1;
wire signed [18-1:0] W_Q2_1_5_2;reg signed [18-1:0] reg_W_Q2_1_5_2=1128;reg stb_W_Q2_1_5_2;assign W_Q2_1_5_2=reg_W_Q2_1_5_2;
wire signed [18-1:0] W_Q2_1_5_3;reg signed [18-1:0] reg_W_Q2_1_5_3=259316;reg stb_W_Q2_1_5_3;assign W_Q2_1_5_3=reg_W_Q2_1_5_3;
wire signed [18-1:0] W_Q2_1_6_0;reg signed [18-1:0] reg_W_Q2_1_6_0=796;reg stb_W_Q2_1_6_0;assign W_Q2_1_6_0=reg_W_Q2_1_6_0;
wire signed [18-1:0] W_Q2_1_6_1;reg signed [18-1:0] reg_W_Q2_1_6_1=9162;reg stb_W_Q2_1_6_1;assign W_Q2_1_6_1=reg_W_Q2_1_6_1;
wire signed [18-1:0] W_Q2_1_6_2;reg signed [18-1:0] reg_W_Q2_1_6_2=260588;reg stb_W_Q2_1_6_2;assign W_Q2_1_6_2=reg_W_Q2_1_6_2;
wire signed [18-1:0] W_Q2_1_6_3;reg signed [18-1:0] reg_W_Q2_1_6_3=13399;reg stb_W_Q2_1_6_3;assign W_Q2_1_6_3=reg_W_Q2_1_6_3;
wire signed [18-1:0] W_Q2_1_7_0;reg signed [18-1:0] reg_W_Q2_1_7_0=2316;reg stb_W_Q2_1_7_0;assign W_Q2_1_7_0=reg_W_Q2_1_7_0;
wire signed [18-1:0] W_Q2_1_7_1;reg signed [18-1:0] reg_W_Q2_1_7_1=11726;reg stb_W_Q2_1_7_1;assign W_Q2_1_7_1=reg_W_Q2_1_7_1;
wire signed [18-1:0] W_Q2_1_7_2;reg signed [18-1:0] reg_W_Q2_1_7_2=80;reg stb_W_Q2_1_7_2;assign W_Q2_1_7_2=reg_W_Q2_1_7_2;
wire signed [18-1:0] W_Q2_1_7_3;reg signed [18-1:0] reg_W_Q2_1_7_3=8325;reg stb_W_Q2_1_7_3;assign W_Q2_1_7_3=reg_W_Q2_1_7_3;
wire signed [18-1:0] W_Q2_2_0_0;reg signed [18-1:0] reg_W_Q2_2_0_0=3299;reg stb_W_Q2_2_0_0;assign W_Q2_2_0_0=reg_W_Q2_2_0_0;
wire signed [18-1:0] W_Q2_2_1_0;reg signed [18-1:0] reg_W_Q2_2_1_0=247774;reg stb_W_Q2_2_1_0;assign W_Q2_2_1_0=reg_W_Q2_2_1_0;
wire signed [18-1:0] W_Q2_2_2_0;reg signed [18-1:0] reg_W_Q2_2_2_0=258016;reg stb_W_Q2_2_2_0;assign W_Q2_2_2_0=reg_W_Q2_2_2_0;
wire signed [18-1:0] W_Q2_2_3_0;reg signed [18-1:0] reg_W_Q2_2_3_0=248723;reg stb_W_Q2_2_3_0;assign W_Q2_2_3_0=reg_W_Q2_2_3_0;
wire signed [18-1:0] B_Q2_0_0;reg signed [18-1:0] reg_B_Q2_0_0=262042;reg stb_B_Q2_0_0;assign B_Q2_0_0=reg_B_Q2_0_0;
wire signed [18-1:0] B_Q2_0_1;reg signed [18-1:0] reg_B_Q2_0_1=259230;reg stb_B_Q2_0_1;assign B_Q2_0_1=reg_B_Q2_0_1;
wire signed [18-1:0] B_Q2_0_2;reg signed [18-1:0] reg_B_Q2_0_2=0;reg stb_B_Q2_0_2;assign B_Q2_0_2=reg_B_Q2_0_2;
wire signed [18-1:0] B_Q2_0_3;reg signed [18-1:0] reg_B_Q2_0_3=0;reg stb_B_Q2_0_3;assign B_Q2_0_3=reg_B_Q2_0_3;
wire signed [18-1:0] B_Q2_0_4;reg signed [18-1:0] reg_B_Q2_0_4=0;reg stb_B_Q2_0_4;assign B_Q2_0_4=reg_B_Q2_0_4;
wire signed [18-1:0] B_Q2_0_5;reg signed [18-1:0] reg_B_Q2_0_5=0;reg stb_B_Q2_0_5;assign B_Q2_0_5=reg_B_Q2_0_5;
wire signed [18-1:0] B_Q2_0_6;reg signed [18-1:0] reg_B_Q2_0_6=258988;reg stb_B_Q2_0_6;assign B_Q2_0_6=reg_B_Q2_0_6;
wire signed [18-1:0] B_Q2_0_7;reg signed [18-1:0] reg_B_Q2_0_7=259290;reg stb_B_Q2_0_7;assign B_Q2_0_7=reg_B_Q2_0_7;
wire signed [18-1:0] B_Q2_1_0;reg signed [18-1:0] reg_B_Q2_1_0=262129;reg stb_B_Q2_1_0;assign B_Q2_1_0=reg_B_Q2_1_0;
wire signed [18-1:0] B_Q2_1_1;reg signed [18-1:0] reg_B_Q2_1_1=259931;reg stb_B_Q2_1_1;assign B_Q2_1_1=reg_B_Q2_1_1;
wire signed [18-1:0] B_Q2_1_2;reg signed [18-1:0] reg_B_Q2_1_2=0;reg stb_B_Q2_1_2;assign B_Q2_1_2=reg_B_Q2_1_2;
wire signed [18-1:0] B_Q2_1_3;reg signed [18-1:0] reg_B_Q2_1_3=259739;reg stb_B_Q2_1_3;assign B_Q2_1_3=reg_B_Q2_1_3;
wire signed [18-1:0] B_Q2_2_0;reg signed [18-1:0] reg_B_Q2_2_0=22860;reg stb_B_Q2_2_0;assign B_Q2_2_0=reg_B_Q2_2_0;
wire signed [18-1:0] W_Q3_0_0_0;reg signed [18-1:0] reg_W_Q3_0_0_0=260183;reg stb_W_Q3_0_0_0;assign W_Q3_0_0_0=reg_W_Q3_0_0_0;
wire signed [18-1:0] W_Q3_0_0_1;reg signed [18-1:0] reg_W_Q3_0_0_1=4862;reg stb_W_Q3_0_0_1;assign W_Q3_0_0_1=reg_W_Q3_0_0_1;
wire signed [18-1:0] W_Q3_0_0_2;reg signed [18-1:0] reg_W_Q3_0_0_2=261334;reg stb_W_Q3_0_0_2;assign W_Q3_0_0_2=reg_W_Q3_0_0_2;
wire signed [18-1:0] W_Q3_0_0_3;reg signed [18-1:0] reg_W_Q3_0_0_3=260711;reg stb_W_Q3_0_0_3;assign W_Q3_0_0_3=reg_W_Q3_0_0_3;
wire signed [18-1:0] W_Q3_0_0_4;reg signed [18-1:0] reg_W_Q3_0_0_4=262141;reg stb_W_Q3_0_0_4;assign W_Q3_0_0_4=reg_W_Q3_0_0_4;
wire signed [18-1:0] W_Q3_0_0_5;reg signed [18-1:0] reg_W_Q3_0_0_5=259938;reg stb_W_Q3_0_0_5;assign W_Q3_0_0_5=reg_W_Q3_0_0_5;
wire signed [18-1:0] W_Q3_0_0_6;reg signed [18-1:0] reg_W_Q3_0_0_6=4215;reg stb_W_Q3_0_0_6;assign W_Q3_0_0_6=reg_W_Q3_0_0_6;
wire signed [18-1:0] W_Q3_0_0_7;reg signed [18-1:0] reg_W_Q3_0_0_7=4895;reg stb_W_Q3_0_0_7;assign W_Q3_0_0_7=reg_W_Q3_0_0_7;
wire signed [18-1:0] W_Q3_0_1_0;reg signed [18-1:0] reg_W_Q3_0_1_0=1258;reg stb_W_Q3_0_1_0;assign W_Q3_0_1_0=reg_W_Q3_0_1_0;
wire signed [18-1:0] W_Q3_0_1_1;reg signed [18-1:0] reg_W_Q3_0_1_1=4406;reg stb_W_Q3_0_1_1;assign W_Q3_0_1_1=reg_W_Q3_0_1_1;
wire signed [18-1:0] W_Q3_0_1_2;reg signed [18-1:0] reg_W_Q3_0_1_2=259194;reg stb_W_Q3_0_1_2;assign W_Q3_0_1_2=reg_W_Q3_0_1_2;
wire signed [18-1:0] W_Q3_0_1_3;reg signed [18-1:0] reg_W_Q3_0_1_3=260609;reg stb_W_Q3_0_1_3;assign W_Q3_0_1_3=reg_W_Q3_0_1_3;
wire signed [18-1:0] W_Q3_0_1_4;reg signed [18-1:0] reg_W_Q3_0_1_4=260881;reg stb_W_Q3_0_1_4;assign W_Q3_0_1_4=reg_W_Q3_0_1_4;
wire signed [18-1:0] W_Q3_0_1_5;reg signed [18-1:0] reg_W_Q3_0_1_5=261883;reg stb_W_Q3_0_1_5;assign W_Q3_0_1_5=reg_W_Q3_0_1_5;
wire signed [18-1:0] W_Q3_0_1_6;reg signed [18-1:0] reg_W_Q3_0_1_6=3074;reg stb_W_Q3_0_1_6;assign W_Q3_0_1_6=reg_W_Q3_0_1_6;
wire signed [18-1:0] W_Q3_0_1_7;reg signed [18-1:0] reg_W_Q3_0_1_7=2106;reg stb_W_Q3_0_1_7;assign W_Q3_0_1_7=reg_W_Q3_0_1_7;
wire signed [18-1:0] W_Q3_1_0_0;reg signed [18-1:0] reg_W_Q3_1_0_0=260105;reg stb_W_Q3_1_0_0;assign W_Q3_1_0_0=reg_W_Q3_1_0_0;
wire signed [18-1:0] W_Q3_1_0_1;reg signed [18-1:0] reg_W_Q3_1_0_1=261076;reg stb_W_Q3_1_0_1;assign W_Q3_1_0_1=reg_W_Q3_1_0_1;
wire signed [18-1:0] W_Q3_1_0_2;reg signed [18-1:0] reg_W_Q3_1_0_2=1240;reg stb_W_Q3_1_0_2;assign W_Q3_1_0_2=reg_W_Q3_1_0_2;
wire signed [18-1:0] W_Q3_1_0_3;reg signed [18-1:0] reg_W_Q3_1_0_3=2377;reg stb_W_Q3_1_0_3;assign W_Q3_1_0_3=reg_W_Q3_1_0_3;
wire signed [18-1:0] W_Q3_1_1_0;reg signed [18-1:0] reg_W_Q3_1_1_0=260362;reg stb_W_Q3_1_1_0;assign W_Q3_1_1_0=reg_W_Q3_1_1_0;
wire signed [18-1:0] W_Q3_1_1_1;reg signed [18-1:0] reg_W_Q3_1_1_1=6050;reg stb_W_Q3_1_1_1;assign W_Q3_1_1_1=reg_W_Q3_1_1_1;
wire signed [18-1:0] W_Q3_1_1_2;reg signed [18-1:0] reg_W_Q3_1_1_2=261792;reg stb_W_Q3_1_1_2;assign W_Q3_1_1_2=reg_W_Q3_1_1_2;
wire signed [18-1:0] W_Q3_1_1_3;reg signed [18-1:0] reg_W_Q3_1_1_3=7072;reg stb_W_Q3_1_1_3;assign W_Q3_1_1_3=reg_W_Q3_1_1_3;
wire signed [18-1:0] W_Q3_1_2_0;reg signed [18-1:0] reg_W_Q3_1_2_0=261219;reg stb_W_Q3_1_2_0;assign W_Q3_1_2_0=reg_W_Q3_1_2_0;
wire signed [18-1:0] W_Q3_1_2_1;reg signed [18-1:0] reg_W_Q3_1_2_1=261083;reg stb_W_Q3_1_2_1;assign W_Q3_1_2_1=reg_W_Q3_1_2_1;
wire signed [18-1:0] W_Q3_1_2_2;reg signed [18-1:0] reg_W_Q3_1_2_2=231;reg stb_W_Q3_1_2_2;assign W_Q3_1_2_2=reg_W_Q3_1_2_2;
wire signed [18-1:0] W_Q3_1_2_3;reg signed [18-1:0] reg_W_Q3_1_2_3=2514;reg stb_W_Q3_1_2_3;assign W_Q3_1_2_3=reg_W_Q3_1_2_3;
wire signed [18-1:0] W_Q3_1_3_0;reg signed [18-1:0] reg_W_Q3_1_3_0=1992;reg stb_W_Q3_1_3_0;assign W_Q3_1_3_0=reg_W_Q3_1_3_0;
wire signed [18-1:0] W_Q3_1_3_1;reg signed [18-1:0] reg_W_Q3_1_3_1=2883;reg stb_W_Q3_1_3_1;assign W_Q3_1_3_1=reg_W_Q3_1_3_1;
wire signed [18-1:0] W_Q3_1_3_2;reg signed [18-1:0] reg_W_Q3_1_3_2=260124;reg stb_W_Q3_1_3_2;assign W_Q3_1_3_2=reg_W_Q3_1_3_2;
wire signed [18-1:0] W_Q3_1_3_3;reg signed [18-1:0] reg_W_Q3_1_3_3=260161;reg stb_W_Q3_1_3_3;assign W_Q3_1_3_3=reg_W_Q3_1_3_3;
wire signed [18-1:0] W_Q3_1_4_0;reg signed [18-1:0] reg_W_Q3_1_4_0=260317;reg stb_W_Q3_1_4_0;assign W_Q3_1_4_0=reg_W_Q3_1_4_0;
wire signed [18-1:0] W_Q3_1_4_1;reg signed [18-1:0] reg_W_Q3_1_4_1=259731;reg stb_W_Q3_1_4_1;assign W_Q3_1_4_1=reg_W_Q3_1_4_1;
wire signed [18-1:0] W_Q3_1_4_2;reg signed [18-1:0] reg_W_Q3_1_4_2=261824;reg stb_W_Q3_1_4_2;assign W_Q3_1_4_2=reg_W_Q3_1_4_2;
wire signed [18-1:0] W_Q3_1_4_3;reg signed [18-1:0] reg_W_Q3_1_4_3=261593;reg stb_W_Q3_1_4_3;assign W_Q3_1_4_3=reg_W_Q3_1_4_3;
wire signed [18-1:0] W_Q3_1_5_0;reg signed [18-1:0] reg_W_Q3_1_5_0=2757;reg stb_W_Q3_1_5_0;assign W_Q3_1_5_0=reg_W_Q3_1_5_0;
wire signed [18-1:0] W_Q3_1_5_1;reg signed [18-1:0] reg_W_Q3_1_5_1=261239;reg stb_W_Q3_1_5_1;assign W_Q3_1_5_1=reg_W_Q3_1_5_1;
wire signed [18-1:0] W_Q3_1_5_2;reg signed [18-1:0] reg_W_Q3_1_5_2=1128;reg stb_W_Q3_1_5_2;assign W_Q3_1_5_2=reg_W_Q3_1_5_2;
wire signed [18-1:0] W_Q3_1_5_3;reg signed [18-1:0] reg_W_Q3_1_5_3=259316;reg stb_W_Q3_1_5_3;assign W_Q3_1_5_3=reg_W_Q3_1_5_3;
wire signed [18-1:0] W_Q3_1_6_0;reg signed [18-1:0] reg_W_Q3_1_6_0=796;reg stb_W_Q3_1_6_0;assign W_Q3_1_6_0=reg_W_Q3_1_6_0;
wire signed [18-1:0] W_Q3_1_6_1;reg signed [18-1:0] reg_W_Q3_1_6_1=9162;reg stb_W_Q3_1_6_1;assign W_Q3_1_6_1=reg_W_Q3_1_6_1;
wire signed [18-1:0] W_Q3_1_6_2;reg signed [18-1:0] reg_W_Q3_1_6_2=260588;reg stb_W_Q3_1_6_2;assign W_Q3_1_6_2=reg_W_Q3_1_6_2;
wire signed [18-1:0] W_Q3_1_6_3;reg signed [18-1:0] reg_W_Q3_1_6_3=13399;reg stb_W_Q3_1_6_3;assign W_Q3_1_6_3=reg_W_Q3_1_6_3;
wire signed [18-1:0] W_Q3_1_7_0;reg signed [18-1:0] reg_W_Q3_1_7_0=2316;reg stb_W_Q3_1_7_0;assign W_Q3_1_7_0=reg_W_Q3_1_7_0;
wire signed [18-1:0] W_Q3_1_7_1;reg signed [18-1:0] reg_W_Q3_1_7_1=11726;reg stb_W_Q3_1_7_1;assign W_Q3_1_7_1=reg_W_Q3_1_7_1;
wire signed [18-1:0] W_Q3_1_7_2;reg signed [18-1:0] reg_W_Q3_1_7_2=80;reg stb_W_Q3_1_7_2;assign W_Q3_1_7_2=reg_W_Q3_1_7_2;
wire signed [18-1:0] W_Q3_1_7_3;reg signed [18-1:0] reg_W_Q3_1_7_3=8325;reg stb_W_Q3_1_7_3;assign W_Q3_1_7_3=reg_W_Q3_1_7_3;
wire signed [18-1:0] W_Q3_2_0_0;reg signed [18-1:0] reg_W_Q3_2_0_0=3299;reg stb_W_Q3_2_0_0;assign W_Q3_2_0_0=reg_W_Q3_2_0_0;
wire signed [18-1:0] W_Q3_2_1_0;reg signed [18-1:0] reg_W_Q3_2_1_0=247774;reg stb_W_Q3_2_1_0;assign W_Q3_2_1_0=reg_W_Q3_2_1_0;
wire signed [18-1:0] W_Q3_2_2_0;reg signed [18-1:0] reg_W_Q3_2_2_0=258016;reg stb_W_Q3_2_2_0;assign W_Q3_2_2_0=reg_W_Q3_2_2_0;
wire signed [18-1:0] W_Q3_2_3_0;reg signed [18-1:0] reg_W_Q3_2_3_0=248723;reg stb_W_Q3_2_3_0;assign W_Q3_2_3_0=reg_W_Q3_2_3_0;
wire signed [18-1:0] B_Q3_0_0;reg signed [18-1:0] reg_B_Q3_0_0=262042;reg stb_B_Q3_0_0;assign B_Q3_0_0=reg_B_Q3_0_0;
wire signed [18-1:0] B_Q3_0_1;reg signed [18-1:0] reg_B_Q3_0_1=259230;reg stb_B_Q3_0_1;assign B_Q3_0_1=reg_B_Q3_0_1;
wire signed [18-1:0] B_Q3_0_2;reg signed [18-1:0] reg_B_Q3_0_2=0;reg stb_B_Q3_0_2;assign B_Q3_0_2=reg_B_Q3_0_2;
wire signed [18-1:0] B_Q3_0_3;reg signed [18-1:0] reg_B_Q3_0_3=0;reg stb_B_Q3_0_3;assign B_Q3_0_3=reg_B_Q3_0_3;
wire signed [18-1:0] B_Q3_0_4;reg signed [18-1:0] reg_B_Q3_0_4=0;reg stb_B_Q3_0_4;assign B_Q3_0_4=reg_B_Q3_0_4;
wire signed [18-1:0] B_Q3_0_5;reg signed [18-1:0] reg_B_Q3_0_5=0;reg stb_B_Q3_0_5;assign B_Q3_0_5=reg_B_Q3_0_5;
wire signed [18-1:0] B_Q3_0_6;reg signed [18-1:0] reg_B_Q3_0_6=258988;reg stb_B_Q3_0_6;assign B_Q3_0_6=reg_B_Q3_0_6;
wire signed [18-1:0] B_Q3_0_7;reg signed [18-1:0] reg_B_Q3_0_7=259290;reg stb_B_Q3_0_7;assign B_Q3_0_7=reg_B_Q3_0_7;
wire signed [18-1:0] B_Q3_1_0;reg signed [18-1:0] reg_B_Q3_1_0=262129;reg stb_B_Q3_1_0;assign B_Q3_1_0=reg_B_Q3_1_0;
wire signed [18-1:0] B_Q3_1_1;reg signed [18-1:0] reg_B_Q3_1_1=259931;reg stb_B_Q3_1_1;assign B_Q3_1_1=reg_B_Q3_1_1;
wire signed [18-1:0] B_Q3_1_2;reg signed [18-1:0] reg_B_Q3_1_2=0;reg stb_B_Q3_1_2;assign B_Q3_1_2=reg_B_Q3_1_2;
wire signed [18-1:0] B_Q3_1_3;reg signed [18-1:0] reg_B_Q3_1_3=259739;reg stb_B_Q3_1_3;assign B_Q3_1_3=reg_B_Q3_1_3;
wire signed [18-1:0] B_Q3_2_0;reg signed [18-1:0] reg_B_Q3_2_0=22860;reg stb_B_Q3_2_0;assign B_Q3_2_0=reg_B_Q3_2_0;
wire signed [18-1:0] W_Q4_0_0_0;reg signed [18-1:0] reg_W_Q4_0_0_0=260183;reg stb_W_Q4_0_0_0;assign W_Q4_0_0_0=reg_W_Q4_0_0_0;
wire signed [18-1:0] W_Q4_0_0_1;reg signed [18-1:0] reg_W_Q4_0_0_1=4862;reg stb_W_Q4_0_0_1;assign W_Q4_0_0_1=reg_W_Q4_0_0_1;
wire signed [18-1:0] W_Q4_0_0_2;reg signed [18-1:0] reg_W_Q4_0_0_2=261334;reg stb_W_Q4_0_0_2;assign W_Q4_0_0_2=reg_W_Q4_0_0_2;
wire signed [18-1:0] W_Q4_0_0_3;reg signed [18-1:0] reg_W_Q4_0_0_3=260711;reg stb_W_Q4_0_0_3;assign W_Q4_0_0_3=reg_W_Q4_0_0_3;
wire signed [18-1:0] W_Q4_0_0_4;reg signed [18-1:0] reg_W_Q4_0_0_4=262141;reg stb_W_Q4_0_0_4;assign W_Q4_0_0_4=reg_W_Q4_0_0_4;
wire signed [18-1:0] W_Q4_0_0_5;reg signed [18-1:0] reg_W_Q4_0_0_5=259938;reg stb_W_Q4_0_0_5;assign W_Q4_0_0_5=reg_W_Q4_0_0_5;
wire signed [18-1:0] W_Q4_0_0_6;reg signed [18-1:0] reg_W_Q4_0_0_6=4215;reg stb_W_Q4_0_0_6;assign W_Q4_0_0_6=reg_W_Q4_0_0_6;
wire signed [18-1:0] W_Q4_0_0_7;reg signed [18-1:0] reg_W_Q4_0_0_7=4895;reg stb_W_Q4_0_0_7;assign W_Q4_0_0_7=reg_W_Q4_0_0_7;
wire signed [18-1:0] W_Q4_0_1_0;reg signed [18-1:0] reg_W_Q4_0_1_0=1258;reg stb_W_Q4_0_1_0;assign W_Q4_0_1_0=reg_W_Q4_0_1_0;
wire signed [18-1:0] W_Q4_0_1_1;reg signed [18-1:0] reg_W_Q4_0_1_1=4406;reg stb_W_Q4_0_1_1;assign W_Q4_0_1_1=reg_W_Q4_0_1_1;
wire signed [18-1:0] W_Q4_0_1_2;reg signed [18-1:0] reg_W_Q4_0_1_2=259194;reg stb_W_Q4_0_1_2;assign W_Q4_0_1_2=reg_W_Q4_0_1_2;
wire signed [18-1:0] W_Q4_0_1_3;reg signed [18-1:0] reg_W_Q4_0_1_3=260609;reg stb_W_Q4_0_1_3;assign W_Q4_0_1_3=reg_W_Q4_0_1_3;
wire signed [18-1:0] W_Q4_0_1_4;reg signed [18-1:0] reg_W_Q4_0_1_4=260881;reg stb_W_Q4_0_1_4;assign W_Q4_0_1_4=reg_W_Q4_0_1_4;
wire signed [18-1:0] W_Q4_0_1_5;reg signed [18-1:0] reg_W_Q4_0_1_5=261883;reg stb_W_Q4_0_1_5;assign W_Q4_0_1_5=reg_W_Q4_0_1_5;
wire signed [18-1:0] W_Q4_0_1_6;reg signed [18-1:0] reg_W_Q4_0_1_6=3074;reg stb_W_Q4_0_1_6;assign W_Q4_0_1_6=reg_W_Q4_0_1_6;
wire signed [18-1:0] W_Q4_0_1_7;reg signed [18-1:0] reg_W_Q4_0_1_7=2106;reg stb_W_Q4_0_1_7;assign W_Q4_0_1_7=reg_W_Q4_0_1_7;
wire signed [18-1:0] W_Q4_1_0_0;reg signed [18-1:0] reg_W_Q4_1_0_0=260105;reg stb_W_Q4_1_0_0;assign W_Q4_1_0_0=reg_W_Q4_1_0_0;
wire signed [18-1:0] W_Q4_1_0_1;reg signed [18-1:0] reg_W_Q4_1_0_1=261076;reg stb_W_Q4_1_0_1;assign W_Q4_1_0_1=reg_W_Q4_1_0_1;
wire signed [18-1:0] W_Q4_1_0_2;reg signed [18-1:0] reg_W_Q4_1_0_2=1240;reg stb_W_Q4_1_0_2;assign W_Q4_1_0_2=reg_W_Q4_1_0_2;
wire signed [18-1:0] W_Q4_1_0_3;reg signed [18-1:0] reg_W_Q4_1_0_3=2377;reg stb_W_Q4_1_0_3;assign W_Q4_1_0_3=reg_W_Q4_1_0_3;
wire signed [18-1:0] W_Q4_1_1_0;reg signed [18-1:0] reg_W_Q4_1_1_0=260362;reg stb_W_Q4_1_1_0;assign W_Q4_1_1_0=reg_W_Q4_1_1_0;
wire signed [18-1:0] W_Q4_1_1_1;reg signed [18-1:0] reg_W_Q4_1_1_1=6050;reg stb_W_Q4_1_1_1;assign W_Q4_1_1_1=reg_W_Q4_1_1_1;
wire signed [18-1:0] W_Q4_1_1_2;reg signed [18-1:0] reg_W_Q4_1_1_2=261792;reg stb_W_Q4_1_1_2;assign W_Q4_1_1_2=reg_W_Q4_1_1_2;
wire signed [18-1:0] W_Q4_1_1_3;reg signed [18-1:0] reg_W_Q4_1_1_3=7072;reg stb_W_Q4_1_1_3;assign W_Q4_1_1_3=reg_W_Q4_1_1_3;
wire signed [18-1:0] W_Q4_1_2_0;reg signed [18-1:0] reg_W_Q4_1_2_0=261219;reg stb_W_Q4_1_2_0;assign W_Q4_1_2_0=reg_W_Q4_1_2_0;
wire signed [18-1:0] W_Q4_1_2_1;reg signed [18-1:0] reg_W_Q4_1_2_1=261083;reg stb_W_Q4_1_2_1;assign W_Q4_1_2_1=reg_W_Q4_1_2_1;
wire signed [18-1:0] W_Q4_1_2_2;reg signed [18-1:0] reg_W_Q4_1_2_2=231;reg stb_W_Q4_1_2_2;assign W_Q4_1_2_2=reg_W_Q4_1_2_2;
wire signed [18-1:0] W_Q4_1_2_3;reg signed [18-1:0] reg_W_Q4_1_2_3=2514;reg stb_W_Q4_1_2_3;assign W_Q4_1_2_3=reg_W_Q4_1_2_3;
wire signed [18-1:0] W_Q4_1_3_0;reg signed [18-1:0] reg_W_Q4_1_3_0=1992;reg stb_W_Q4_1_3_0;assign W_Q4_1_3_0=reg_W_Q4_1_3_0;
wire signed [18-1:0] W_Q4_1_3_1;reg signed [18-1:0] reg_W_Q4_1_3_1=2883;reg stb_W_Q4_1_3_1;assign W_Q4_1_3_1=reg_W_Q4_1_3_1;
wire signed [18-1:0] W_Q4_1_3_2;reg signed [18-1:0] reg_W_Q4_1_3_2=260124;reg stb_W_Q4_1_3_2;assign W_Q4_1_3_2=reg_W_Q4_1_3_2;
wire signed [18-1:0] W_Q4_1_3_3;reg signed [18-1:0] reg_W_Q4_1_3_3=260161;reg stb_W_Q4_1_3_3;assign W_Q4_1_3_3=reg_W_Q4_1_3_3;
wire signed [18-1:0] W_Q4_1_4_0;reg signed [18-1:0] reg_W_Q4_1_4_0=260317;reg stb_W_Q4_1_4_0;assign W_Q4_1_4_0=reg_W_Q4_1_4_0;
wire signed [18-1:0] W_Q4_1_4_1;reg signed [18-1:0] reg_W_Q4_1_4_1=259731;reg stb_W_Q4_1_4_1;assign W_Q4_1_4_1=reg_W_Q4_1_4_1;
wire signed [18-1:0] W_Q4_1_4_2;reg signed [18-1:0] reg_W_Q4_1_4_2=261824;reg stb_W_Q4_1_4_2;assign W_Q4_1_4_2=reg_W_Q4_1_4_2;
wire signed [18-1:0] W_Q4_1_4_3;reg signed [18-1:0] reg_W_Q4_1_4_3=261593;reg stb_W_Q4_1_4_3;assign W_Q4_1_4_3=reg_W_Q4_1_4_3;
wire signed [18-1:0] W_Q4_1_5_0;reg signed [18-1:0] reg_W_Q4_1_5_0=2757;reg stb_W_Q4_1_5_0;assign W_Q4_1_5_0=reg_W_Q4_1_5_0;
wire signed [18-1:0] W_Q4_1_5_1;reg signed [18-1:0] reg_W_Q4_1_5_1=261239;reg stb_W_Q4_1_5_1;assign W_Q4_1_5_1=reg_W_Q4_1_5_1;
wire signed [18-1:0] W_Q4_1_5_2;reg signed [18-1:0] reg_W_Q4_1_5_2=1128;reg stb_W_Q4_1_5_2;assign W_Q4_1_5_2=reg_W_Q4_1_5_2;
wire signed [18-1:0] W_Q4_1_5_3;reg signed [18-1:0] reg_W_Q4_1_5_3=259316;reg stb_W_Q4_1_5_3;assign W_Q4_1_5_3=reg_W_Q4_1_5_3;
wire signed [18-1:0] W_Q4_1_6_0;reg signed [18-1:0] reg_W_Q4_1_6_0=796;reg stb_W_Q4_1_6_0;assign W_Q4_1_6_0=reg_W_Q4_1_6_0;
wire signed [18-1:0] W_Q4_1_6_1;reg signed [18-1:0] reg_W_Q4_1_6_1=9162;reg stb_W_Q4_1_6_1;assign W_Q4_1_6_1=reg_W_Q4_1_6_1;
wire signed [18-1:0] W_Q4_1_6_2;reg signed [18-1:0] reg_W_Q4_1_6_2=260588;reg stb_W_Q4_1_6_2;assign W_Q4_1_6_2=reg_W_Q4_1_6_2;
wire signed [18-1:0] W_Q4_1_6_3;reg signed [18-1:0] reg_W_Q4_1_6_3=13399;reg stb_W_Q4_1_6_3;assign W_Q4_1_6_3=reg_W_Q4_1_6_3;
wire signed [18-1:0] W_Q4_1_7_0;reg signed [18-1:0] reg_W_Q4_1_7_0=2316;reg stb_W_Q4_1_7_0;assign W_Q4_1_7_0=reg_W_Q4_1_7_0;
wire signed [18-1:0] W_Q4_1_7_1;reg signed [18-1:0] reg_W_Q4_1_7_1=11726;reg stb_W_Q4_1_7_1;assign W_Q4_1_7_1=reg_W_Q4_1_7_1;
wire signed [18-1:0] W_Q4_1_7_2;reg signed [18-1:0] reg_W_Q4_1_7_2=80;reg stb_W_Q4_1_7_2;assign W_Q4_1_7_2=reg_W_Q4_1_7_2;
wire signed [18-1:0] W_Q4_1_7_3;reg signed [18-1:0] reg_W_Q4_1_7_3=8325;reg stb_W_Q4_1_7_3;assign W_Q4_1_7_3=reg_W_Q4_1_7_3;
wire signed [18-1:0] W_Q4_2_0_0;reg signed [18-1:0] reg_W_Q4_2_0_0=3299;reg stb_W_Q4_2_0_0;assign W_Q4_2_0_0=reg_W_Q4_2_0_0;
wire signed [18-1:0] W_Q4_2_1_0;reg signed [18-1:0] reg_W_Q4_2_1_0=247774;reg stb_W_Q4_2_1_0;assign W_Q4_2_1_0=reg_W_Q4_2_1_0;
wire signed [18-1:0] W_Q4_2_2_0;reg signed [18-1:0] reg_W_Q4_2_2_0=258016;reg stb_W_Q4_2_2_0;assign W_Q4_2_2_0=reg_W_Q4_2_2_0;
wire signed [18-1:0] W_Q4_2_3_0;reg signed [18-1:0] reg_W_Q4_2_3_0=248723;reg stb_W_Q4_2_3_0;assign W_Q4_2_3_0=reg_W_Q4_2_3_0;
wire signed [18-1:0] B_Q4_0_0;reg signed [18-1:0] reg_B_Q4_0_0=262042;reg stb_B_Q4_0_0;assign B_Q4_0_0=reg_B_Q4_0_0;
wire signed [18-1:0] B_Q4_0_1;reg signed [18-1:0] reg_B_Q4_0_1=259230;reg stb_B_Q4_0_1;assign B_Q4_0_1=reg_B_Q4_0_1;
wire signed [18-1:0] B_Q4_0_2;reg signed [18-1:0] reg_B_Q4_0_2=0;reg stb_B_Q4_0_2;assign B_Q4_0_2=reg_B_Q4_0_2;
wire signed [18-1:0] B_Q4_0_3;reg signed [18-1:0] reg_B_Q4_0_3=0;reg stb_B_Q4_0_3;assign B_Q4_0_3=reg_B_Q4_0_3;
wire signed [18-1:0] B_Q4_0_4;reg signed [18-1:0] reg_B_Q4_0_4=0;reg stb_B_Q4_0_4;assign B_Q4_0_4=reg_B_Q4_0_4;
wire signed [18-1:0] B_Q4_0_5;reg signed [18-1:0] reg_B_Q4_0_5=0;reg stb_B_Q4_0_5;assign B_Q4_0_5=reg_B_Q4_0_5;
wire signed [18-1:0] B_Q4_0_6;reg signed [18-1:0] reg_B_Q4_0_6=258988;reg stb_B_Q4_0_6;assign B_Q4_0_6=reg_B_Q4_0_6;
wire signed [18-1:0] B_Q4_0_7;reg signed [18-1:0] reg_B_Q4_0_7=259290;reg stb_B_Q4_0_7;assign B_Q4_0_7=reg_B_Q4_0_7;
wire signed [18-1:0] B_Q4_1_0;reg signed [18-1:0] reg_B_Q4_1_0=262129;reg stb_B_Q4_1_0;assign B_Q4_1_0=reg_B_Q4_1_0;
wire signed [18-1:0] B_Q4_1_1;reg signed [18-1:0] reg_B_Q4_1_1=259931;reg stb_B_Q4_1_1;assign B_Q4_1_1=reg_B_Q4_1_1;
wire signed [18-1:0] B_Q4_1_2;reg signed [18-1:0] reg_B_Q4_1_2=0;reg stb_B_Q4_1_2;assign B_Q4_1_2=reg_B_Q4_1_2;
wire signed [18-1:0] B_Q4_1_3;reg signed [18-1:0] reg_B_Q4_1_3=259739;reg stb_B_Q4_1_3;assign B_Q4_1_3=reg_B_Q4_1_3;
wire signed [18-1:0] B_Q4_2_0;reg signed [18-1:0] reg_B_Q4_2_0=22860;reg stb_B_Q4_2_0;assign B_Q4_2_0=reg_B_Q4_2_0;
wire signed [18-1:0] W_Q5_0_0_0;reg signed [18-1:0] reg_W_Q5_0_0_0=260183;reg stb_W_Q5_0_0_0;assign W_Q5_0_0_0=reg_W_Q5_0_0_0;
wire signed [18-1:0] W_Q5_0_0_1;reg signed [18-1:0] reg_W_Q5_0_0_1=4862;reg stb_W_Q5_0_0_1;assign W_Q5_0_0_1=reg_W_Q5_0_0_1;
wire signed [18-1:0] W_Q5_0_0_2;reg signed [18-1:0] reg_W_Q5_0_0_2=261334;reg stb_W_Q5_0_0_2;assign W_Q5_0_0_2=reg_W_Q5_0_0_2;
wire signed [18-1:0] W_Q5_0_0_3;reg signed [18-1:0] reg_W_Q5_0_0_3=260711;reg stb_W_Q5_0_0_3;assign W_Q5_0_0_3=reg_W_Q5_0_0_3;
wire signed [18-1:0] W_Q5_0_0_4;reg signed [18-1:0] reg_W_Q5_0_0_4=262141;reg stb_W_Q5_0_0_4;assign W_Q5_0_0_4=reg_W_Q5_0_0_4;
wire signed [18-1:0] W_Q5_0_0_5;reg signed [18-1:0] reg_W_Q5_0_0_5=259938;reg stb_W_Q5_0_0_5;assign W_Q5_0_0_5=reg_W_Q5_0_0_5;
wire signed [18-1:0] W_Q5_0_0_6;reg signed [18-1:0] reg_W_Q5_0_0_6=4215;reg stb_W_Q5_0_0_6;assign W_Q5_0_0_6=reg_W_Q5_0_0_6;
wire signed [18-1:0] W_Q5_0_0_7;reg signed [18-1:0] reg_W_Q5_0_0_7=4895;reg stb_W_Q5_0_0_7;assign W_Q5_0_0_7=reg_W_Q5_0_0_7;
wire signed [18-1:0] W_Q5_0_1_0;reg signed [18-1:0] reg_W_Q5_0_1_0=1258;reg stb_W_Q5_0_1_0;assign W_Q5_0_1_0=reg_W_Q5_0_1_0;
wire signed [18-1:0] W_Q5_0_1_1;reg signed [18-1:0] reg_W_Q5_0_1_1=4406;reg stb_W_Q5_0_1_1;assign W_Q5_0_1_1=reg_W_Q5_0_1_1;
wire signed [18-1:0] W_Q5_0_1_2;reg signed [18-1:0] reg_W_Q5_0_1_2=259194;reg stb_W_Q5_0_1_2;assign W_Q5_0_1_2=reg_W_Q5_0_1_2;
wire signed [18-1:0] W_Q5_0_1_3;reg signed [18-1:0] reg_W_Q5_0_1_3=260609;reg stb_W_Q5_0_1_3;assign W_Q5_0_1_3=reg_W_Q5_0_1_3;
wire signed [18-1:0] W_Q5_0_1_4;reg signed [18-1:0] reg_W_Q5_0_1_4=260881;reg stb_W_Q5_0_1_4;assign W_Q5_0_1_4=reg_W_Q5_0_1_4;
wire signed [18-1:0] W_Q5_0_1_5;reg signed [18-1:0] reg_W_Q5_0_1_5=261883;reg stb_W_Q5_0_1_5;assign W_Q5_0_1_5=reg_W_Q5_0_1_5;
wire signed [18-1:0] W_Q5_0_1_6;reg signed [18-1:0] reg_W_Q5_0_1_6=3074;reg stb_W_Q5_0_1_6;assign W_Q5_0_1_6=reg_W_Q5_0_1_6;
wire signed [18-1:0] W_Q5_0_1_7;reg signed [18-1:0] reg_W_Q5_0_1_7=2106;reg stb_W_Q5_0_1_7;assign W_Q5_0_1_7=reg_W_Q5_0_1_7;
wire signed [18-1:0] W_Q5_1_0_0;reg signed [18-1:0] reg_W_Q5_1_0_0=260105;reg stb_W_Q5_1_0_0;assign W_Q5_1_0_0=reg_W_Q5_1_0_0;
wire signed [18-1:0] W_Q5_1_0_1;reg signed [18-1:0] reg_W_Q5_1_0_1=261076;reg stb_W_Q5_1_0_1;assign W_Q5_1_0_1=reg_W_Q5_1_0_1;
wire signed [18-1:0] W_Q5_1_0_2;reg signed [18-1:0] reg_W_Q5_1_0_2=1240;reg stb_W_Q5_1_0_2;assign W_Q5_1_0_2=reg_W_Q5_1_0_2;
wire signed [18-1:0] W_Q5_1_0_3;reg signed [18-1:0] reg_W_Q5_1_0_3=2377;reg stb_W_Q5_1_0_3;assign W_Q5_1_0_3=reg_W_Q5_1_0_3;
wire signed [18-1:0] W_Q5_1_1_0;reg signed [18-1:0] reg_W_Q5_1_1_0=260362;reg stb_W_Q5_1_1_0;assign W_Q5_1_1_0=reg_W_Q5_1_1_0;
wire signed [18-1:0] W_Q5_1_1_1;reg signed [18-1:0] reg_W_Q5_1_1_1=6050;reg stb_W_Q5_1_1_1;assign W_Q5_1_1_1=reg_W_Q5_1_1_1;
wire signed [18-1:0] W_Q5_1_1_2;reg signed [18-1:0] reg_W_Q5_1_1_2=261792;reg stb_W_Q5_1_1_2;assign W_Q5_1_1_2=reg_W_Q5_1_1_2;
wire signed [18-1:0] W_Q5_1_1_3;reg signed [18-1:0] reg_W_Q5_1_1_3=7072;reg stb_W_Q5_1_1_3;assign W_Q5_1_1_3=reg_W_Q5_1_1_3;
wire signed [18-1:0] W_Q5_1_2_0;reg signed [18-1:0] reg_W_Q5_1_2_0=261219;reg stb_W_Q5_1_2_0;assign W_Q5_1_2_0=reg_W_Q5_1_2_0;
wire signed [18-1:0] W_Q5_1_2_1;reg signed [18-1:0] reg_W_Q5_1_2_1=261083;reg stb_W_Q5_1_2_1;assign W_Q5_1_2_1=reg_W_Q5_1_2_1;
wire signed [18-1:0] W_Q5_1_2_2;reg signed [18-1:0] reg_W_Q5_1_2_2=231;reg stb_W_Q5_1_2_2;assign W_Q5_1_2_2=reg_W_Q5_1_2_2;
wire signed [18-1:0] W_Q5_1_2_3;reg signed [18-1:0] reg_W_Q5_1_2_3=2514;reg stb_W_Q5_1_2_3;assign W_Q5_1_2_3=reg_W_Q5_1_2_3;
wire signed [18-1:0] W_Q5_1_3_0;reg signed [18-1:0] reg_W_Q5_1_3_0=1992;reg stb_W_Q5_1_3_0;assign W_Q5_1_3_0=reg_W_Q5_1_3_0;
wire signed [18-1:0] W_Q5_1_3_1;reg signed [18-1:0] reg_W_Q5_1_3_1=2883;reg stb_W_Q5_1_3_1;assign W_Q5_1_3_1=reg_W_Q5_1_3_1;
wire signed [18-1:0] W_Q5_1_3_2;reg signed [18-1:0] reg_W_Q5_1_3_2=260124;reg stb_W_Q5_1_3_2;assign W_Q5_1_3_2=reg_W_Q5_1_3_2;
wire signed [18-1:0] W_Q5_1_3_3;reg signed [18-1:0] reg_W_Q5_1_3_3=260161;reg stb_W_Q5_1_3_3;assign W_Q5_1_3_3=reg_W_Q5_1_3_3;
wire signed [18-1:0] W_Q5_1_4_0;reg signed [18-1:0] reg_W_Q5_1_4_0=260317;reg stb_W_Q5_1_4_0;assign W_Q5_1_4_0=reg_W_Q5_1_4_0;
wire signed [18-1:0] W_Q5_1_4_1;reg signed [18-1:0] reg_W_Q5_1_4_1=259731;reg stb_W_Q5_1_4_1;assign W_Q5_1_4_1=reg_W_Q5_1_4_1;
wire signed [18-1:0] W_Q5_1_4_2;reg signed [18-1:0] reg_W_Q5_1_4_2=261824;reg stb_W_Q5_1_4_2;assign W_Q5_1_4_2=reg_W_Q5_1_4_2;
wire signed [18-1:0] W_Q5_1_4_3;reg signed [18-1:0] reg_W_Q5_1_4_3=261593;reg stb_W_Q5_1_4_3;assign W_Q5_1_4_3=reg_W_Q5_1_4_3;
wire signed [18-1:0] W_Q5_1_5_0;reg signed [18-1:0] reg_W_Q5_1_5_0=2757;reg stb_W_Q5_1_5_0;assign W_Q5_1_5_0=reg_W_Q5_1_5_0;
wire signed [18-1:0] W_Q5_1_5_1;reg signed [18-1:0] reg_W_Q5_1_5_1=261239;reg stb_W_Q5_1_5_1;assign W_Q5_1_5_1=reg_W_Q5_1_5_1;
wire signed [18-1:0] W_Q5_1_5_2;reg signed [18-1:0] reg_W_Q5_1_5_2=1128;reg stb_W_Q5_1_5_2;assign W_Q5_1_5_2=reg_W_Q5_1_5_2;
wire signed [18-1:0] W_Q5_1_5_3;reg signed [18-1:0] reg_W_Q5_1_5_3=259316;reg stb_W_Q5_1_5_3;assign W_Q5_1_5_3=reg_W_Q5_1_5_3;
wire signed [18-1:0] W_Q5_1_6_0;reg signed [18-1:0] reg_W_Q5_1_6_0=796;reg stb_W_Q5_1_6_0;assign W_Q5_1_6_0=reg_W_Q5_1_6_0;
wire signed [18-1:0] W_Q5_1_6_1;reg signed [18-1:0] reg_W_Q5_1_6_1=9162;reg stb_W_Q5_1_6_1;assign W_Q5_1_6_1=reg_W_Q5_1_6_1;
wire signed [18-1:0] W_Q5_1_6_2;reg signed [18-1:0] reg_W_Q5_1_6_2=260588;reg stb_W_Q5_1_6_2;assign W_Q5_1_6_2=reg_W_Q5_1_6_2;
wire signed [18-1:0] W_Q5_1_6_3;reg signed [18-1:0] reg_W_Q5_1_6_3=13399;reg stb_W_Q5_1_6_3;assign W_Q5_1_6_3=reg_W_Q5_1_6_3;
wire signed [18-1:0] W_Q5_1_7_0;reg signed [18-1:0] reg_W_Q5_1_7_0=2316;reg stb_W_Q5_1_7_0;assign W_Q5_1_7_0=reg_W_Q5_1_7_0;
wire signed [18-1:0] W_Q5_1_7_1;reg signed [18-1:0] reg_W_Q5_1_7_1=11726;reg stb_W_Q5_1_7_1;assign W_Q5_1_7_1=reg_W_Q5_1_7_1;
wire signed [18-1:0] W_Q5_1_7_2;reg signed [18-1:0] reg_W_Q5_1_7_2=80;reg stb_W_Q5_1_7_2;assign W_Q5_1_7_2=reg_W_Q5_1_7_2;
wire signed [18-1:0] W_Q5_1_7_3;reg signed [18-1:0] reg_W_Q5_1_7_3=8325;reg stb_W_Q5_1_7_3;assign W_Q5_1_7_3=reg_W_Q5_1_7_3;
wire signed [18-1:0] W_Q5_2_0_0;reg signed [18-1:0] reg_W_Q5_2_0_0=3299;reg stb_W_Q5_2_0_0;assign W_Q5_2_0_0=reg_W_Q5_2_0_0;
wire signed [18-1:0] W_Q5_2_1_0;reg signed [18-1:0] reg_W_Q5_2_1_0=247774;reg stb_W_Q5_2_1_0;assign W_Q5_2_1_0=reg_W_Q5_2_1_0;
wire signed [18-1:0] W_Q5_2_2_0;reg signed [18-1:0] reg_W_Q5_2_2_0=258016;reg stb_W_Q5_2_2_0;assign W_Q5_2_2_0=reg_W_Q5_2_2_0;
wire signed [18-1:0] W_Q5_2_3_0;reg signed [18-1:0] reg_W_Q5_2_3_0=248723;reg stb_W_Q5_2_3_0;assign W_Q5_2_3_0=reg_W_Q5_2_3_0;
wire signed [18-1:0] B_Q5_0_0;reg signed [18-1:0] reg_B_Q5_0_0=262042;reg stb_B_Q5_0_0;assign B_Q5_0_0=reg_B_Q5_0_0;
wire signed [18-1:0] B_Q5_0_1;reg signed [18-1:0] reg_B_Q5_0_1=259230;reg stb_B_Q5_0_1;assign B_Q5_0_1=reg_B_Q5_0_1;
wire signed [18-1:0] B_Q5_0_2;reg signed [18-1:0] reg_B_Q5_0_2=0;reg stb_B_Q5_0_2;assign B_Q5_0_2=reg_B_Q5_0_2;
wire signed [18-1:0] B_Q5_0_3;reg signed [18-1:0] reg_B_Q5_0_3=0;reg stb_B_Q5_0_3;assign B_Q5_0_3=reg_B_Q5_0_3;
wire signed [18-1:0] B_Q5_0_4;reg signed [18-1:0] reg_B_Q5_0_4=0;reg stb_B_Q5_0_4;assign B_Q5_0_4=reg_B_Q5_0_4;
wire signed [18-1:0] B_Q5_0_5;reg signed [18-1:0] reg_B_Q5_0_5=0;reg stb_B_Q5_0_5;assign B_Q5_0_5=reg_B_Q5_0_5;
wire signed [18-1:0] B_Q5_0_6;reg signed [18-1:0] reg_B_Q5_0_6=258988;reg stb_B_Q5_0_6;assign B_Q5_0_6=reg_B_Q5_0_6;
wire signed [18-1:0] B_Q5_0_7;reg signed [18-1:0] reg_B_Q5_0_7=259290;reg stb_B_Q5_0_7;assign B_Q5_0_7=reg_B_Q5_0_7;
wire signed [18-1:0] B_Q5_1_0;reg signed [18-1:0] reg_B_Q5_1_0=262129;reg stb_B_Q5_1_0;assign B_Q5_1_0=reg_B_Q5_1_0;
wire signed [18-1:0] B_Q5_1_1;reg signed [18-1:0] reg_B_Q5_1_1=259931;reg stb_B_Q5_1_1;assign B_Q5_1_1=reg_B_Q5_1_1;
wire signed [18-1:0] B_Q5_1_2;reg signed [18-1:0] reg_B_Q5_1_2=0;reg stb_B_Q5_1_2;assign B_Q5_1_2=reg_B_Q5_1_2;
wire signed [18-1:0] B_Q5_1_3;reg signed [18-1:0] reg_B_Q5_1_3=259739;reg stb_B_Q5_1_3;assign B_Q5_1_3=reg_B_Q5_1_3;
wire signed [18-1:0] B_Q5_2_0;reg signed [18-1:0] reg_B_Q5_2_0=22860;reg stb_B_Q5_2_0;assign B_Q5_2_0=reg_B_Q5_2_0;
wire signed [18-1:0] W_Q6_0_0_0;reg signed [18-1:0] reg_W_Q6_0_0_0=260183;reg stb_W_Q6_0_0_0;assign W_Q6_0_0_0=reg_W_Q6_0_0_0;
wire signed [18-1:0] W_Q6_0_0_1;reg signed [18-1:0] reg_W_Q6_0_0_1=4862;reg stb_W_Q6_0_0_1;assign W_Q6_0_0_1=reg_W_Q6_0_0_1;
wire signed [18-1:0] W_Q6_0_0_2;reg signed [18-1:0] reg_W_Q6_0_0_2=261334;reg stb_W_Q6_0_0_2;assign W_Q6_0_0_2=reg_W_Q6_0_0_2;
wire signed [18-1:0] W_Q6_0_0_3;reg signed [18-1:0] reg_W_Q6_0_0_3=260711;reg stb_W_Q6_0_0_3;assign W_Q6_0_0_3=reg_W_Q6_0_0_3;
wire signed [18-1:0] W_Q6_0_0_4;reg signed [18-1:0] reg_W_Q6_0_0_4=262141;reg stb_W_Q6_0_0_4;assign W_Q6_0_0_4=reg_W_Q6_0_0_4;
wire signed [18-1:0] W_Q6_0_0_5;reg signed [18-1:0] reg_W_Q6_0_0_5=259938;reg stb_W_Q6_0_0_5;assign W_Q6_0_0_5=reg_W_Q6_0_0_5;
wire signed [18-1:0] W_Q6_0_0_6;reg signed [18-1:0] reg_W_Q6_0_0_6=4215;reg stb_W_Q6_0_0_6;assign W_Q6_0_0_6=reg_W_Q6_0_0_6;
wire signed [18-1:0] W_Q6_0_0_7;reg signed [18-1:0] reg_W_Q6_0_0_7=4895;reg stb_W_Q6_0_0_7;assign W_Q6_0_0_7=reg_W_Q6_0_0_7;
wire signed [18-1:0] W_Q6_0_1_0;reg signed [18-1:0] reg_W_Q6_0_1_0=1258;reg stb_W_Q6_0_1_0;assign W_Q6_0_1_0=reg_W_Q6_0_1_0;
wire signed [18-1:0] W_Q6_0_1_1;reg signed [18-1:0] reg_W_Q6_0_1_1=4406;reg stb_W_Q6_0_1_1;assign W_Q6_0_1_1=reg_W_Q6_0_1_1;
wire signed [18-1:0] W_Q6_0_1_2;reg signed [18-1:0] reg_W_Q6_0_1_2=259194;reg stb_W_Q6_0_1_2;assign W_Q6_0_1_2=reg_W_Q6_0_1_2;
wire signed [18-1:0] W_Q6_0_1_3;reg signed [18-1:0] reg_W_Q6_0_1_3=260609;reg stb_W_Q6_0_1_3;assign W_Q6_0_1_3=reg_W_Q6_0_1_3;
wire signed [18-1:0] W_Q6_0_1_4;reg signed [18-1:0] reg_W_Q6_0_1_4=260881;reg stb_W_Q6_0_1_4;assign W_Q6_0_1_4=reg_W_Q6_0_1_4;
wire signed [18-1:0] W_Q6_0_1_5;reg signed [18-1:0] reg_W_Q6_0_1_5=261883;reg stb_W_Q6_0_1_5;assign W_Q6_0_1_5=reg_W_Q6_0_1_5;
wire signed [18-1:0] W_Q6_0_1_6;reg signed [18-1:0] reg_W_Q6_0_1_6=3074;reg stb_W_Q6_0_1_6;assign W_Q6_0_1_6=reg_W_Q6_0_1_6;
wire signed [18-1:0] W_Q6_0_1_7;reg signed [18-1:0] reg_W_Q6_0_1_7=2106;reg stb_W_Q6_0_1_7;assign W_Q6_0_1_7=reg_W_Q6_0_1_7;
wire signed [18-1:0] W_Q6_1_0_0;reg signed [18-1:0] reg_W_Q6_1_0_0=260105;reg stb_W_Q6_1_0_0;assign W_Q6_1_0_0=reg_W_Q6_1_0_0;
wire signed [18-1:0] W_Q6_1_0_1;reg signed [18-1:0] reg_W_Q6_1_0_1=261076;reg stb_W_Q6_1_0_1;assign W_Q6_1_0_1=reg_W_Q6_1_0_1;
wire signed [18-1:0] W_Q6_1_0_2;reg signed [18-1:0] reg_W_Q6_1_0_2=1240;reg stb_W_Q6_1_0_2;assign W_Q6_1_0_2=reg_W_Q6_1_0_2;
wire signed [18-1:0] W_Q6_1_0_3;reg signed [18-1:0] reg_W_Q6_1_0_3=2377;reg stb_W_Q6_1_0_3;assign W_Q6_1_0_3=reg_W_Q6_1_0_3;
wire signed [18-1:0] W_Q6_1_1_0;reg signed [18-1:0] reg_W_Q6_1_1_0=260362;reg stb_W_Q6_1_1_0;assign W_Q6_1_1_0=reg_W_Q6_1_1_0;
wire signed [18-1:0] W_Q6_1_1_1;reg signed [18-1:0] reg_W_Q6_1_1_1=6050;reg stb_W_Q6_1_1_1;assign W_Q6_1_1_1=reg_W_Q6_1_1_1;
wire signed [18-1:0] W_Q6_1_1_2;reg signed [18-1:0] reg_W_Q6_1_1_2=261792;reg stb_W_Q6_1_1_2;assign W_Q6_1_1_2=reg_W_Q6_1_1_2;
wire signed [18-1:0] W_Q6_1_1_3;reg signed [18-1:0] reg_W_Q6_1_1_3=7072;reg stb_W_Q6_1_1_3;assign W_Q6_1_1_3=reg_W_Q6_1_1_3;
wire signed [18-1:0] W_Q6_1_2_0;reg signed [18-1:0] reg_W_Q6_1_2_0=261219;reg stb_W_Q6_1_2_0;assign W_Q6_1_2_0=reg_W_Q6_1_2_0;
wire signed [18-1:0] W_Q6_1_2_1;reg signed [18-1:0] reg_W_Q6_1_2_1=261083;reg stb_W_Q6_1_2_1;assign W_Q6_1_2_1=reg_W_Q6_1_2_1;
wire signed [18-1:0] W_Q6_1_2_2;reg signed [18-1:0] reg_W_Q6_1_2_2=231;reg stb_W_Q6_1_2_2;assign W_Q6_1_2_2=reg_W_Q6_1_2_2;
wire signed [18-1:0] W_Q6_1_2_3;reg signed [18-1:0] reg_W_Q6_1_2_3=2514;reg stb_W_Q6_1_2_3;assign W_Q6_1_2_3=reg_W_Q6_1_2_3;
wire signed [18-1:0] W_Q6_1_3_0;reg signed [18-1:0] reg_W_Q6_1_3_0=1992;reg stb_W_Q6_1_3_0;assign W_Q6_1_3_0=reg_W_Q6_1_3_0;
wire signed [18-1:0] W_Q6_1_3_1;reg signed [18-1:0] reg_W_Q6_1_3_1=2883;reg stb_W_Q6_1_3_1;assign W_Q6_1_3_1=reg_W_Q6_1_3_1;
wire signed [18-1:0] W_Q6_1_3_2;reg signed [18-1:0] reg_W_Q6_1_3_2=260124;reg stb_W_Q6_1_3_2;assign W_Q6_1_3_2=reg_W_Q6_1_3_2;
wire signed [18-1:0] W_Q6_1_3_3;reg signed [18-1:0] reg_W_Q6_1_3_3=260161;reg stb_W_Q6_1_3_3;assign W_Q6_1_3_3=reg_W_Q6_1_3_3;
wire signed [18-1:0] W_Q6_1_4_0;reg signed [18-1:0] reg_W_Q6_1_4_0=260317;reg stb_W_Q6_1_4_0;assign W_Q6_1_4_0=reg_W_Q6_1_4_0;
wire signed [18-1:0] W_Q6_1_4_1;reg signed [18-1:0] reg_W_Q6_1_4_1=259731;reg stb_W_Q6_1_4_1;assign W_Q6_1_4_1=reg_W_Q6_1_4_1;
wire signed [18-1:0] W_Q6_1_4_2;reg signed [18-1:0] reg_W_Q6_1_4_2=261824;reg stb_W_Q6_1_4_2;assign W_Q6_1_4_2=reg_W_Q6_1_4_2;
wire signed [18-1:0] W_Q6_1_4_3;reg signed [18-1:0] reg_W_Q6_1_4_3=261593;reg stb_W_Q6_1_4_3;assign W_Q6_1_4_3=reg_W_Q6_1_4_3;
wire signed [18-1:0] W_Q6_1_5_0;reg signed [18-1:0] reg_W_Q6_1_5_0=2757;reg stb_W_Q6_1_5_0;assign W_Q6_1_5_0=reg_W_Q6_1_5_0;
wire signed [18-1:0] W_Q6_1_5_1;reg signed [18-1:0] reg_W_Q6_1_5_1=261239;reg stb_W_Q6_1_5_1;assign W_Q6_1_5_1=reg_W_Q6_1_5_1;
wire signed [18-1:0] W_Q6_1_5_2;reg signed [18-1:0] reg_W_Q6_1_5_2=1128;reg stb_W_Q6_1_5_2;assign W_Q6_1_5_2=reg_W_Q6_1_5_2;
wire signed [18-1:0] W_Q6_1_5_3;reg signed [18-1:0] reg_W_Q6_1_5_3=259316;reg stb_W_Q6_1_5_3;assign W_Q6_1_5_3=reg_W_Q6_1_5_3;
wire signed [18-1:0] W_Q6_1_6_0;reg signed [18-1:0] reg_W_Q6_1_6_0=796;reg stb_W_Q6_1_6_0;assign W_Q6_1_6_0=reg_W_Q6_1_6_0;
wire signed [18-1:0] W_Q6_1_6_1;reg signed [18-1:0] reg_W_Q6_1_6_1=9162;reg stb_W_Q6_1_6_1;assign W_Q6_1_6_1=reg_W_Q6_1_6_1;
wire signed [18-1:0] W_Q6_1_6_2;reg signed [18-1:0] reg_W_Q6_1_6_2=260588;reg stb_W_Q6_1_6_2;assign W_Q6_1_6_2=reg_W_Q6_1_6_2;
wire signed [18-1:0] W_Q6_1_6_3;reg signed [18-1:0] reg_W_Q6_1_6_3=13399;reg stb_W_Q6_1_6_3;assign W_Q6_1_6_3=reg_W_Q6_1_6_3;
wire signed [18-1:0] W_Q6_1_7_0;reg signed [18-1:0] reg_W_Q6_1_7_0=2316;reg stb_W_Q6_1_7_0;assign W_Q6_1_7_0=reg_W_Q6_1_7_0;
wire signed [18-1:0] W_Q6_1_7_1;reg signed [18-1:0] reg_W_Q6_1_7_1=11726;reg stb_W_Q6_1_7_1;assign W_Q6_1_7_1=reg_W_Q6_1_7_1;
wire signed [18-1:0] W_Q6_1_7_2;reg signed [18-1:0] reg_W_Q6_1_7_2=80;reg stb_W_Q6_1_7_2;assign W_Q6_1_7_2=reg_W_Q6_1_7_2;
wire signed [18-1:0] W_Q6_1_7_3;reg signed [18-1:0] reg_W_Q6_1_7_3=8325;reg stb_W_Q6_1_7_3;assign W_Q6_1_7_3=reg_W_Q6_1_7_3;
wire signed [18-1:0] W_Q6_2_0_0;reg signed [18-1:0] reg_W_Q6_2_0_0=3299;reg stb_W_Q6_2_0_0;assign W_Q6_2_0_0=reg_W_Q6_2_0_0;
wire signed [18-1:0] W_Q6_2_1_0;reg signed [18-1:0] reg_W_Q6_2_1_0=247774;reg stb_W_Q6_2_1_0;assign W_Q6_2_1_0=reg_W_Q6_2_1_0;
wire signed [18-1:0] W_Q6_2_2_0;reg signed [18-1:0] reg_W_Q6_2_2_0=258016;reg stb_W_Q6_2_2_0;assign W_Q6_2_2_0=reg_W_Q6_2_2_0;
wire signed [18-1:0] W_Q6_2_3_0;reg signed [18-1:0] reg_W_Q6_2_3_0=248723;reg stb_W_Q6_2_3_0;assign W_Q6_2_3_0=reg_W_Q6_2_3_0;
wire signed [18-1:0] B_Q6_0_0;reg signed [18-1:0] reg_B_Q6_0_0=262042;reg stb_B_Q6_0_0;assign B_Q6_0_0=reg_B_Q6_0_0;
wire signed [18-1:0] B_Q6_0_1;reg signed [18-1:0] reg_B_Q6_0_1=259230;reg stb_B_Q6_0_1;assign B_Q6_0_1=reg_B_Q6_0_1;
wire signed [18-1:0] B_Q6_0_2;reg signed [18-1:0] reg_B_Q6_0_2=0;reg stb_B_Q6_0_2;assign B_Q6_0_2=reg_B_Q6_0_2;
wire signed [18-1:0] B_Q6_0_3;reg signed [18-1:0] reg_B_Q6_0_3=0;reg stb_B_Q6_0_3;assign B_Q6_0_3=reg_B_Q6_0_3;
wire signed [18-1:0] B_Q6_0_4;reg signed [18-1:0] reg_B_Q6_0_4=0;reg stb_B_Q6_0_4;assign B_Q6_0_4=reg_B_Q6_0_4;
wire signed [18-1:0] B_Q6_0_5;reg signed [18-1:0] reg_B_Q6_0_5=0;reg stb_B_Q6_0_5;assign B_Q6_0_5=reg_B_Q6_0_5;
wire signed [18-1:0] B_Q6_0_6;reg signed [18-1:0] reg_B_Q6_0_6=258988;reg stb_B_Q6_0_6;assign B_Q6_0_6=reg_B_Q6_0_6;
wire signed [18-1:0] B_Q6_0_7;reg signed [18-1:0] reg_B_Q6_0_7=259290;reg stb_B_Q6_0_7;assign B_Q6_0_7=reg_B_Q6_0_7;
wire signed [18-1:0] B_Q6_1_0;reg signed [18-1:0] reg_B_Q6_1_0=262129;reg stb_B_Q6_1_0;assign B_Q6_1_0=reg_B_Q6_1_0;
wire signed [18-1:0] B_Q6_1_1;reg signed [18-1:0] reg_B_Q6_1_1=259931;reg stb_B_Q6_1_1;assign B_Q6_1_1=reg_B_Q6_1_1;
wire signed [18-1:0] B_Q6_1_2;reg signed [18-1:0] reg_B_Q6_1_2=0;reg stb_B_Q6_1_2;assign B_Q6_1_2=reg_B_Q6_1_2;
wire signed [18-1:0] B_Q6_1_3;reg signed [18-1:0] reg_B_Q6_1_3=259739;reg stb_B_Q6_1_3;assign B_Q6_1_3=reg_B_Q6_1_3;
wire signed [18-1:0] B_Q6_2_0;reg signed [18-1:0] reg_B_Q6_2_0=22860;reg stb_B_Q6_2_0;assign B_Q6_2_0=reg_B_Q6_2_0;
wire signed [18-1:0] W_Q7_0_0_0;reg signed [18-1:0] reg_W_Q7_0_0_0=260183;reg stb_W_Q7_0_0_0;assign W_Q7_0_0_0=reg_W_Q7_0_0_0;
wire signed [18-1:0] W_Q7_0_0_1;reg signed [18-1:0] reg_W_Q7_0_0_1=4862;reg stb_W_Q7_0_0_1;assign W_Q7_0_0_1=reg_W_Q7_0_0_1;
wire signed [18-1:0] W_Q7_0_0_2;reg signed [18-1:0] reg_W_Q7_0_0_2=261334;reg stb_W_Q7_0_0_2;assign W_Q7_0_0_2=reg_W_Q7_0_0_2;
wire signed [18-1:0] W_Q7_0_0_3;reg signed [18-1:0] reg_W_Q7_0_0_3=260711;reg stb_W_Q7_0_0_3;assign W_Q7_0_0_3=reg_W_Q7_0_0_3;
wire signed [18-1:0] W_Q7_0_0_4;reg signed [18-1:0] reg_W_Q7_0_0_4=262141;reg stb_W_Q7_0_0_4;assign W_Q7_0_0_4=reg_W_Q7_0_0_4;
wire signed [18-1:0] W_Q7_0_0_5;reg signed [18-1:0] reg_W_Q7_0_0_5=259938;reg stb_W_Q7_0_0_5;assign W_Q7_0_0_5=reg_W_Q7_0_0_5;
wire signed [18-1:0] W_Q7_0_0_6;reg signed [18-1:0] reg_W_Q7_0_0_6=4215;reg stb_W_Q7_0_0_6;assign W_Q7_0_0_6=reg_W_Q7_0_0_6;
wire signed [18-1:0] W_Q7_0_0_7;reg signed [18-1:0] reg_W_Q7_0_0_7=4895;reg stb_W_Q7_0_0_7;assign W_Q7_0_0_7=reg_W_Q7_0_0_7;
wire signed [18-1:0] W_Q7_0_1_0;reg signed [18-1:0] reg_W_Q7_0_1_0=1258;reg stb_W_Q7_0_1_0;assign W_Q7_0_1_0=reg_W_Q7_0_1_0;
wire signed [18-1:0] W_Q7_0_1_1;reg signed [18-1:0] reg_W_Q7_0_1_1=4406;reg stb_W_Q7_0_1_1;assign W_Q7_0_1_1=reg_W_Q7_0_1_1;
wire signed [18-1:0] W_Q7_0_1_2;reg signed [18-1:0] reg_W_Q7_0_1_2=259194;reg stb_W_Q7_0_1_2;assign W_Q7_0_1_2=reg_W_Q7_0_1_2;
wire signed [18-1:0] W_Q7_0_1_3;reg signed [18-1:0] reg_W_Q7_0_1_3=260609;reg stb_W_Q7_0_1_3;assign W_Q7_0_1_3=reg_W_Q7_0_1_3;
wire signed [18-1:0] W_Q7_0_1_4;reg signed [18-1:0] reg_W_Q7_0_1_4=260881;reg stb_W_Q7_0_1_4;assign W_Q7_0_1_4=reg_W_Q7_0_1_4;
wire signed [18-1:0] W_Q7_0_1_5;reg signed [18-1:0] reg_W_Q7_0_1_5=261883;reg stb_W_Q7_0_1_5;assign W_Q7_0_1_5=reg_W_Q7_0_1_5;
wire signed [18-1:0] W_Q7_0_1_6;reg signed [18-1:0] reg_W_Q7_0_1_6=3074;reg stb_W_Q7_0_1_6;assign W_Q7_0_1_6=reg_W_Q7_0_1_6;
wire signed [18-1:0] W_Q7_0_1_7;reg signed [18-1:0] reg_W_Q7_0_1_7=2106;reg stb_W_Q7_0_1_7;assign W_Q7_0_1_7=reg_W_Q7_0_1_7;
wire signed [18-1:0] W_Q7_1_0_0;reg signed [18-1:0] reg_W_Q7_1_0_0=260105;reg stb_W_Q7_1_0_0;assign W_Q7_1_0_0=reg_W_Q7_1_0_0;
wire signed [18-1:0] W_Q7_1_0_1;reg signed [18-1:0] reg_W_Q7_1_0_1=261076;reg stb_W_Q7_1_0_1;assign W_Q7_1_0_1=reg_W_Q7_1_0_1;
wire signed [18-1:0] W_Q7_1_0_2;reg signed [18-1:0] reg_W_Q7_1_0_2=1240;reg stb_W_Q7_1_0_2;assign W_Q7_1_0_2=reg_W_Q7_1_0_2;
wire signed [18-1:0] W_Q7_1_0_3;reg signed [18-1:0] reg_W_Q7_1_0_3=2377;reg stb_W_Q7_1_0_3;assign W_Q7_1_0_3=reg_W_Q7_1_0_3;
wire signed [18-1:0] W_Q7_1_1_0;reg signed [18-1:0] reg_W_Q7_1_1_0=260362;reg stb_W_Q7_1_1_0;assign W_Q7_1_1_0=reg_W_Q7_1_1_0;
wire signed [18-1:0] W_Q7_1_1_1;reg signed [18-1:0] reg_W_Q7_1_1_1=6050;reg stb_W_Q7_1_1_1;assign W_Q7_1_1_1=reg_W_Q7_1_1_1;
wire signed [18-1:0] W_Q7_1_1_2;reg signed [18-1:0] reg_W_Q7_1_1_2=261792;reg stb_W_Q7_1_1_2;assign W_Q7_1_1_2=reg_W_Q7_1_1_2;
wire signed [18-1:0] W_Q7_1_1_3;reg signed [18-1:0] reg_W_Q7_1_1_3=7072;reg stb_W_Q7_1_1_3;assign W_Q7_1_1_3=reg_W_Q7_1_1_3;
wire signed [18-1:0] W_Q7_1_2_0;reg signed [18-1:0] reg_W_Q7_1_2_0=261219;reg stb_W_Q7_1_2_0;assign W_Q7_1_2_0=reg_W_Q7_1_2_0;
wire signed [18-1:0] W_Q7_1_2_1;reg signed [18-1:0] reg_W_Q7_1_2_1=261083;reg stb_W_Q7_1_2_1;assign W_Q7_1_2_1=reg_W_Q7_1_2_1;
wire signed [18-1:0] W_Q7_1_2_2;reg signed [18-1:0] reg_W_Q7_1_2_2=231;reg stb_W_Q7_1_2_2;assign W_Q7_1_2_2=reg_W_Q7_1_2_2;
wire signed [18-1:0] W_Q7_1_2_3;reg signed [18-1:0] reg_W_Q7_1_2_3=2514;reg stb_W_Q7_1_2_3;assign W_Q7_1_2_3=reg_W_Q7_1_2_3;
wire signed [18-1:0] W_Q7_1_3_0;reg signed [18-1:0] reg_W_Q7_1_3_0=1992;reg stb_W_Q7_1_3_0;assign W_Q7_1_3_0=reg_W_Q7_1_3_0;
wire signed [18-1:0] W_Q7_1_3_1;reg signed [18-1:0] reg_W_Q7_1_3_1=2883;reg stb_W_Q7_1_3_1;assign W_Q7_1_3_1=reg_W_Q7_1_3_1;
wire signed [18-1:0] W_Q7_1_3_2;reg signed [18-1:0] reg_W_Q7_1_3_2=260124;reg stb_W_Q7_1_3_2;assign W_Q7_1_3_2=reg_W_Q7_1_3_2;
wire signed [18-1:0] W_Q7_1_3_3;reg signed [18-1:0] reg_W_Q7_1_3_3=260161;reg stb_W_Q7_1_3_3;assign W_Q7_1_3_3=reg_W_Q7_1_3_3;
wire signed [18-1:0] W_Q7_1_4_0;reg signed [18-1:0] reg_W_Q7_1_4_0=260317;reg stb_W_Q7_1_4_0;assign W_Q7_1_4_0=reg_W_Q7_1_4_0;
wire signed [18-1:0] W_Q7_1_4_1;reg signed [18-1:0] reg_W_Q7_1_4_1=259731;reg stb_W_Q7_1_4_1;assign W_Q7_1_4_1=reg_W_Q7_1_4_1;
wire signed [18-1:0] W_Q7_1_4_2;reg signed [18-1:0] reg_W_Q7_1_4_2=261824;reg stb_W_Q7_1_4_2;assign W_Q7_1_4_2=reg_W_Q7_1_4_2;
wire signed [18-1:0] W_Q7_1_4_3;reg signed [18-1:0] reg_W_Q7_1_4_3=261593;reg stb_W_Q7_1_4_3;assign W_Q7_1_4_3=reg_W_Q7_1_4_3;
wire signed [18-1:0] W_Q7_1_5_0;reg signed [18-1:0] reg_W_Q7_1_5_0=2757;reg stb_W_Q7_1_5_0;assign W_Q7_1_5_0=reg_W_Q7_1_5_0;
wire signed [18-1:0] W_Q7_1_5_1;reg signed [18-1:0] reg_W_Q7_1_5_1=261239;reg stb_W_Q7_1_5_1;assign W_Q7_1_5_1=reg_W_Q7_1_5_1;
wire signed [18-1:0] W_Q7_1_5_2;reg signed [18-1:0] reg_W_Q7_1_5_2=1128;reg stb_W_Q7_1_5_2;assign W_Q7_1_5_2=reg_W_Q7_1_5_2;
wire signed [18-1:0] W_Q7_1_5_3;reg signed [18-1:0] reg_W_Q7_1_5_3=259316;reg stb_W_Q7_1_5_3;assign W_Q7_1_5_3=reg_W_Q7_1_5_3;
wire signed [18-1:0] W_Q7_1_6_0;reg signed [18-1:0] reg_W_Q7_1_6_0=796;reg stb_W_Q7_1_6_0;assign W_Q7_1_6_0=reg_W_Q7_1_6_0;
wire signed [18-1:0] W_Q7_1_6_1;reg signed [18-1:0] reg_W_Q7_1_6_1=9162;reg stb_W_Q7_1_6_1;assign W_Q7_1_6_1=reg_W_Q7_1_6_1;
wire signed [18-1:0] W_Q7_1_6_2;reg signed [18-1:0] reg_W_Q7_1_6_2=260588;reg stb_W_Q7_1_6_2;assign W_Q7_1_6_2=reg_W_Q7_1_6_2;
wire signed [18-1:0] W_Q7_1_6_3;reg signed [18-1:0] reg_W_Q7_1_6_3=13399;reg stb_W_Q7_1_6_3;assign W_Q7_1_6_3=reg_W_Q7_1_6_3;
wire signed [18-1:0] W_Q7_1_7_0;reg signed [18-1:0] reg_W_Q7_1_7_0=2316;reg stb_W_Q7_1_7_0;assign W_Q7_1_7_0=reg_W_Q7_1_7_0;
wire signed [18-1:0] W_Q7_1_7_1;reg signed [18-1:0] reg_W_Q7_1_7_1=11726;reg stb_W_Q7_1_7_1;assign W_Q7_1_7_1=reg_W_Q7_1_7_1;
wire signed [18-1:0] W_Q7_1_7_2;reg signed [18-1:0] reg_W_Q7_1_7_2=80;reg stb_W_Q7_1_7_2;assign W_Q7_1_7_2=reg_W_Q7_1_7_2;
wire signed [18-1:0] W_Q7_1_7_3;reg signed [18-1:0] reg_W_Q7_1_7_3=8325;reg stb_W_Q7_1_7_3;assign W_Q7_1_7_3=reg_W_Q7_1_7_3;
wire signed [18-1:0] W_Q7_2_0_0;reg signed [18-1:0] reg_W_Q7_2_0_0=3299;reg stb_W_Q7_2_0_0;assign W_Q7_2_0_0=reg_W_Q7_2_0_0;
wire signed [18-1:0] W_Q7_2_1_0;reg signed [18-1:0] reg_W_Q7_2_1_0=247774;reg stb_W_Q7_2_1_0;assign W_Q7_2_1_0=reg_W_Q7_2_1_0;
wire signed [18-1:0] W_Q7_2_2_0;reg signed [18-1:0] reg_W_Q7_2_2_0=258016;reg stb_W_Q7_2_2_0;assign W_Q7_2_2_0=reg_W_Q7_2_2_0;
wire signed [18-1:0] W_Q7_2_3_0;reg signed [18-1:0] reg_W_Q7_2_3_0=248723;reg stb_W_Q7_2_3_0;assign W_Q7_2_3_0=reg_W_Q7_2_3_0;
wire signed [18-1:0] B_Q7_0_0;reg signed [18-1:0] reg_B_Q7_0_0=262042;reg stb_B_Q7_0_0;assign B_Q7_0_0=reg_B_Q7_0_0;
wire signed [18-1:0] B_Q7_0_1;reg signed [18-1:0] reg_B_Q7_0_1=259230;reg stb_B_Q7_0_1;assign B_Q7_0_1=reg_B_Q7_0_1;
wire signed [18-1:0] B_Q7_0_2;reg signed [18-1:0] reg_B_Q7_0_2=0;reg stb_B_Q7_0_2;assign B_Q7_0_2=reg_B_Q7_0_2;
wire signed [18-1:0] B_Q7_0_3;reg signed [18-1:0] reg_B_Q7_0_3=0;reg stb_B_Q7_0_3;assign B_Q7_0_3=reg_B_Q7_0_3;
wire signed [18-1:0] B_Q7_0_4;reg signed [18-1:0] reg_B_Q7_0_4=0;reg stb_B_Q7_0_4;assign B_Q7_0_4=reg_B_Q7_0_4;
wire signed [18-1:0] B_Q7_0_5;reg signed [18-1:0] reg_B_Q7_0_5=0;reg stb_B_Q7_0_5;assign B_Q7_0_5=reg_B_Q7_0_5;
wire signed [18-1:0] B_Q7_0_6;reg signed [18-1:0] reg_B_Q7_0_6=258988;reg stb_B_Q7_0_6;assign B_Q7_0_6=reg_B_Q7_0_6;
wire signed [18-1:0] B_Q7_0_7;reg signed [18-1:0] reg_B_Q7_0_7=259290;reg stb_B_Q7_0_7;assign B_Q7_0_7=reg_B_Q7_0_7;
wire signed [18-1:0] B_Q7_1_0;reg signed [18-1:0] reg_B_Q7_1_0=262129;reg stb_B_Q7_1_0;assign B_Q7_1_0=reg_B_Q7_1_0;
wire signed [18-1:0] B_Q7_1_1;reg signed [18-1:0] reg_B_Q7_1_1=259931;reg stb_B_Q7_1_1;assign B_Q7_1_1=reg_B_Q7_1_1;
wire signed [18-1:0] B_Q7_1_2;reg signed [18-1:0] reg_B_Q7_1_2=0;reg stb_B_Q7_1_2;assign B_Q7_1_2=reg_B_Q7_1_2;
wire signed [18-1:0] B_Q7_1_3;reg signed [18-1:0] reg_B_Q7_1_3=259739;reg stb_B_Q7_1_3;assign B_Q7_1_3=reg_B_Q7_1_3;
wire signed [18-1:0] B_Q7_2_0;reg signed [18-1:0] reg_B_Q7_2_0=22860;reg stb_B_Q7_2_0;assign B_Q7_2_0=reg_B_Q7_2_0;
wire signed [32-1:0] min_Q0_I;reg signed [32-1:0] reg_min_Q0_I=262143;reg stb_min_Q0_I;assign min_Q0_I=reg_min_Q0_I;
wire signed [32-1:0] min_Q0_Q;reg signed [32-1:0] reg_min_Q0_Q=262143;reg stb_min_Q0_Q;assign min_Q0_Q=reg_min_Q0_Q;
wire signed [32-1:0] min_Q1_I;reg signed [32-1:0] reg_min_Q1_I=262143;reg stb_min_Q1_I;assign min_Q1_I=reg_min_Q1_I;
wire signed [32-1:0] min_Q1_Q;reg signed [32-1:0] reg_min_Q1_Q=262143;reg stb_min_Q1_Q;assign min_Q1_Q=reg_min_Q1_Q;
wire signed [32-1:0] min_Q2_I;reg signed [32-1:0] reg_min_Q2_I=262143;reg stb_min_Q2_I;assign min_Q2_I=reg_min_Q2_I;
wire signed [32-1:0] min_Q2_Q;reg signed [32-1:0] reg_min_Q2_Q=262143;reg stb_min_Q2_Q;assign min_Q2_Q=reg_min_Q2_Q;
wire signed [32-1:0] min_Q3_I;reg signed [32-1:0] reg_min_Q3_I=262143;reg stb_min_Q3_I;assign min_Q3_I=reg_min_Q3_I;
wire signed [32-1:0] min_Q3_Q;reg signed [32-1:0] reg_min_Q3_Q=262143;reg stb_min_Q3_Q;assign min_Q3_Q=reg_min_Q3_Q;
wire signed [32-1:0] min_Q4_I;reg signed [32-1:0] reg_min_Q4_I=262143;reg stb_min_Q4_I;assign min_Q4_I=reg_min_Q4_I;
wire signed [32-1:0] min_Q4_Q;reg signed [32-1:0] reg_min_Q4_Q=262143;reg stb_min_Q4_Q;assign min_Q4_Q=reg_min_Q4_Q;
wire signed [32-1:0] min_Q5_I;reg signed [32-1:0] reg_min_Q5_I=262143;reg stb_min_Q5_I;assign min_Q5_I=reg_min_Q5_I;
wire signed [32-1:0] min_Q5_Q;reg signed [32-1:0] reg_min_Q5_Q=262143;reg stb_min_Q5_Q;assign min_Q5_Q=reg_min_Q5_Q;
wire signed [32-1:0] min_Q6_I;reg signed [32-1:0] reg_min_Q6_I=262143;reg stb_min_Q6_I;assign min_Q6_I=reg_min_Q6_I;
wire signed [32-1:0] min_Q6_Q;reg signed [32-1:0] reg_min_Q6_Q=262143;reg stb_min_Q6_Q;assign min_Q6_Q=reg_min_Q6_Q;
wire signed [32-1:0] min_Q7_I;reg signed [32-1:0] reg_min_Q7_I=262143;reg stb_min_Q7_I;assign min_Q7_I=reg_min_Q7_I;
wire signed [32-1:0] min_Q7_Q;reg signed [32-1:0] reg_min_Q7_Q=262143;reg stb_min_Q7_Q;assign min_Q7_Q=reg_min_Q7_Q;
always @(posedge lb.clk) begin
wdata<=lb.wdata;
waddr<=lb.waddr;
wren<=lb.wren;
stb_resetacc<=(lb.waddr==1)&lb.wren;if (stb_resetacc) reg_resetacc<=wdata[32-1:0];
stb_amp<=(lb.waddr==6)&lb.wren;if (stb_amp) reg_amp<=wdata[32-1:0];
stb_bramsel<=(lb.waddr==7)&lb.wren;if (stb_bramsel) reg_bramsel<=wdata[32-1:0];
stb_coef00<=(lb.waddr==9)&lb.wren;if (stb_coef00) reg_coef00<=wdata[32-1:0];
stb_coef01<=(lb.waddr==10)&lb.wren;if (stb_coef01) reg_coef01<=wdata[32-1:0];
stb_coef02<=(lb.waddr==11)&lb.wren;if (stb_coef02) reg_coef02<=wdata[32-1:0];
stb_coef03<=(lb.waddr==12)&lb.wren;if (stb_coef03) reg_coef03<=wdata[32-1:0];
stb_coef10<=(lb.waddr==13)&lb.wren;if (stb_coef10) reg_coef10<=wdata[32-1:0];
stb_coef11<=(lb.waddr==14)&lb.wren;if (stb_coef11) reg_coef11<=wdata[32-1:0];
stb_coef12<=(lb.waddr==15)&lb.wren;if (stb_coef12) reg_coef12<=wdata[32-1:0];
stb_coef13<=(lb.waddr==16)&lb.wren;if (stb_coef13) reg_coef13<=wdata[32-1:0];
stb_coef20<=(lb.waddr==17)&lb.wren;if (stb_coef20) reg_coef20<=wdata[32-1:0];
stb_coef21<=(lb.waddr==18)&lb.wren;if (stb_coef21) reg_coef21<=wdata[32-1:0];
stb_coef22<=(lb.waddr==19)&lb.wren;if (stb_coef22) reg_coef22<=wdata[32-1:0];
stb_coef23<=(lb.waddr==20)&lb.wren;if (stb_coef23) reg_coef23<=wdata[32-1:0];
stb_coef30<=(lb.waddr==21)&lb.wren;if (stb_coef30) reg_coef30<=wdata[32-1:0];
stb_coef31<=(lb.waddr==22)&lb.wren;if (stb_coef31) reg_coef31<=wdata[32-1:0];
stb_coef32<=(lb.waddr==23)&lb.wren;if (stb_coef32) reg_coef32<=wdata[32-1:0];
stb_coef33<=(lb.waddr==24)&lb.wren;if (stb_coef33) reg_coef33<=wdata[32-1:0];
stb_dacsel<=(lb.waddr==25)&lb.wren;if (stb_dacsel) reg_dacsel<=wdata[32-1:0];
stb_dspreset<=(lb.waddr==26)&lb.wren;if (stb_dspreset) reg_dspreset<=wdata[1-1:0];
stb_nshot<=(lb.waddr==28)&lb.wren;if (stb_nshot) reg_nshot<=wdata[32-1:0];
stb_qdrvfreqsel<=(lb.waddr==29)&lb.wren;if (stb_qdrvfreqsel) reg_qdrvfreqsel<=wdata[32-1:0];
stb_rdlofreqsel<=(lb.waddr==30)&lb.wren;if (stb_rdlofreqsel) reg_rdlofreqsel<=wdata[32-1:0];
stb_rdrvfreqsel<=(lb.waddr==31)&lb.wren;if (stb_rdrvfreqsel) reg_rdrvfreqsel<=wdata[32-1:0];
stb_reset_bram_read<=(lb.waddr==32)&lb.wren;if (stb_reset_bram_read) reg_reset_bram_read<=wdata[32-1:0];
stb_start<=(lb.waddr==34)&lb.wren;if (stb_start) reg_start<=wdata[1-1:0];
stb_test<=(lb.waddr==35)&lb.wren;if (stb_test) reg_test<=wdata[32-1:0];
stb_acqbufreset<=(lb.waddr==37)&lb.wren;if (stb_acqbufreset) reg_acqbufreset<=wdata[1-1:0];
stb_dacmonreset<=(lb.waddr==38)&lb.wren;if (stb_dacmonreset) reg_dacmonreset<=wdata[1-1:0];
stb_decimator<=(lb.waddr==39)&lb.wren;if (stb_decimator) reg_decimator<=wdata[8-1:0];
stb_acqchansel0<=(lb.waddr==40)&lb.wren;if (stb_acqchansel0) reg_acqchansel0<=wdata[5-1:0];
stb_acqchansel1<=(lb.waddr==41)&lb.wren;if (stb_acqchansel1) reg_acqchansel1<=wdata[5-1:0];
stb_dacmonchansel0<=(lb.waddr==42)&lb.wren;if (stb_dacmonchansel0) reg_dacmonchansel0<=wdata[5-1:0];
stb_dacmonchansel1<=(lb.waddr==43)&lb.wren;if (stb_dacmonchansel1) reg_dacmonchansel1<=wdata[5-1:0];
stb_dacmonchansel2<=(lb.waddr==44)&lb.wren;if (stb_dacmonchansel2) reg_dacmonchansel2<=wdata[5-1:0];
stb_dacmonchansel3<=(lb.waddr==45)&lb.wren;if (stb_dacmonchansel3) reg_dacmonchansel3<=wdata[5-1:0];
stb_delayaftertrig<=(lb.waddr==46)&lb.wren;if (stb_delayaftertrig) reg_delayaftertrig<=wdata[16-1:0];
stb_mixbb1sel<=(lb.waddr==47)&lb.wren;if (stb_mixbb1sel) reg_mixbb1sel<=wdata[16-1:0];
stb_mixbb2sel<=(lb.waddr==48)&lb.wren;if (stb_mixbb2sel) reg_mixbb2sel<=wdata[16-1:0];
stb_shift<=(lb.waddr==49)&lb.wren;if (stb_shift) reg_shift<=wdata[5-1:0];
stb_W_Q0_0_0_0<=(lb.waddr==69)&lb.wren;if (stb_W_Q0_0_0_0) reg_W_Q0_0_0_0<=wdata[18-1:0];
stb_W_Q0_0_0_1<=(lb.waddr==70)&lb.wren;if (stb_W_Q0_0_0_1) reg_W_Q0_0_0_1<=wdata[18-1:0];
stb_W_Q0_0_0_2<=(lb.waddr==71)&lb.wren;if (stb_W_Q0_0_0_2) reg_W_Q0_0_0_2<=wdata[18-1:0];
stb_W_Q0_0_0_3<=(lb.waddr==72)&lb.wren;if (stb_W_Q0_0_0_3) reg_W_Q0_0_0_3<=wdata[18-1:0];
stb_W_Q0_0_0_4<=(lb.waddr==73)&lb.wren;if (stb_W_Q0_0_0_4) reg_W_Q0_0_0_4<=wdata[18-1:0];
stb_W_Q0_0_0_5<=(lb.waddr==74)&lb.wren;if (stb_W_Q0_0_0_5) reg_W_Q0_0_0_5<=wdata[18-1:0];
stb_W_Q0_0_0_6<=(lb.waddr==75)&lb.wren;if (stb_W_Q0_0_0_6) reg_W_Q0_0_0_6<=wdata[18-1:0];
stb_W_Q0_0_0_7<=(lb.waddr==76)&lb.wren;if (stb_W_Q0_0_0_7) reg_W_Q0_0_0_7<=wdata[18-1:0];
stb_W_Q0_0_1_0<=(lb.waddr==77)&lb.wren;if (stb_W_Q0_0_1_0) reg_W_Q0_0_1_0<=wdata[18-1:0];
stb_W_Q0_0_1_1<=(lb.waddr==78)&lb.wren;if (stb_W_Q0_0_1_1) reg_W_Q0_0_1_1<=wdata[18-1:0];
stb_W_Q0_0_1_2<=(lb.waddr==79)&lb.wren;if (stb_W_Q0_0_1_2) reg_W_Q0_0_1_2<=wdata[18-1:0];
stb_W_Q0_0_1_3<=(lb.waddr==80)&lb.wren;if (stb_W_Q0_0_1_3) reg_W_Q0_0_1_3<=wdata[18-1:0];
stb_W_Q0_0_1_4<=(lb.waddr==81)&lb.wren;if (stb_W_Q0_0_1_4) reg_W_Q0_0_1_4<=wdata[18-1:0];
stb_W_Q0_0_1_5<=(lb.waddr==82)&lb.wren;if (stb_W_Q0_0_1_5) reg_W_Q0_0_1_5<=wdata[18-1:0];
stb_W_Q0_0_1_6<=(lb.waddr==83)&lb.wren;if (stb_W_Q0_0_1_6) reg_W_Q0_0_1_6<=wdata[18-1:0];
stb_W_Q0_0_1_7<=(lb.waddr==84)&lb.wren;if (stb_W_Q0_0_1_7) reg_W_Q0_0_1_7<=wdata[18-1:0];
stb_W_Q0_1_0_0<=(lb.waddr==85)&lb.wren;if (stb_W_Q0_1_0_0) reg_W_Q0_1_0_0<=wdata[18-1:0];
stb_W_Q0_1_0_1<=(lb.waddr==86)&lb.wren;if (stb_W_Q0_1_0_1) reg_W_Q0_1_0_1<=wdata[18-1:0];
stb_W_Q0_1_0_2<=(lb.waddr==87)&lb.wren;if (stb_W_Q0_1_0_2) reg_W_Q0_1_0_2<=wdata[18-1:0];
stb_W_Q0_1_0_3<=(lb.waddr==88)&lb.wren;if (stb_W_Q0_1_0_3) reg_W_Q0_1_0_3<=wdata[18-1:0];
stb_W_Q0_1_1_0<=(lb.waddr==89)&lb.wren;if (stb_W_Q0_1_1_0) reg_W_Q0_1_1_0<=wdata[18-1:0];
stb_W_Q0_1_1_1<=(lb.waddr==90)&lb.wren;if (stb_W_Q0_1_1_1) reg_W_Q0_1_1_1<=wdata[18-1:0];
stb_W_Q0_1_1_2<=(lb.waddr==91)&lb.wren;if (stb_W_Q0_1_1_2) reg_W_Q0_1_1_2<=wdata[18-1:0];
stb_W_Q0_1_1_3<=(lb.waddr==92)&lb.wren;if (stb_W_Q0_1_1_3) reg_W_Q0_1_1_3<=wdata[18-1:0];
stb_W_Q0_1_2_0<=(lb.waddr==93)&lb.wren;if (stb_W_Q0_1_2_0) reg_W_Q0_1_2_0<=wdata[18-1:0];
stb_W_Q0_1_2_1<=(lb.waddr==94)&lb.wren;if (stb_W_Q0_1_2_1) reg_W_Q0_1_2_1<=wdata[18-1:0];
stb_W_Q0_1_2_2<=(lb.waddr==95)&lb.wren;if (stb_W_Q0_1_2_2) reg_W_Q0_1_2_2<=wdata[18-1:0];
stb_W_Q0_1_2_3<=(lb.waddr==96)&lb.wren;if (stb_W_Q0_1_2_3) reg_W_Q0_1_2_3<=wdata[18-1:0];
stb_W_Q0_1_3_0<=(lb.waddr==97)&lb.wren;if (stb_W_Q0_1_3_0) reg_W_Q0_1_3_0<=wdata[18-1:0];
stb_W_Q0_1_3_1<=(lb.waddr==98)&lb.wren;if (stb_W_Q0_1_3_1) reg_W_Q0_1_3_1<=wdata[18-1:0];
stb_W_Q0_1_3_2<=(lb.waddr==99)&lb.wren;if (stb_W_Q0_1_3_2) reg_W_Q0_1_3_2<=wdata[18-1:0];
stb_W_Q0_1_3_3<=(lb.waddr==100)&lb.wren;if (stb_W_Q0_1_3_3) reg_W_Q0_1_3_3<=wdata[18-1:0];
stb_W_Q0_1_4_0<=(lb.waddr==101)&lb.wren;if (stb_W_Q0_1_4_0) reg_W_Q0_1_4_0<=wdata[18-1:0];
stb_W_Q0_1_4_1<=(lb.waddr==102)&lb.wren;if (stb_W_Q0_1_4_1) reg_W_Q0_1_4_1<=wdata[18-1:0];
stb_W_Q0_1_4_2<=(lb.waddr==103)&lb.wren;if (stb_W_Q0_1_4_2) reg_W_Q0_1_4_2<=wdata[18-1:0];
stb_W_Q0_1_4_3<=(lb.waddr==104)&lb.wren;if (stb_W_Q0_1_4_3) reg_W_Q0_1_4_3<=wdata[18-1:0];
stb_W_Q0_1_5_0<=(lb.waddr==105)&lb.wren;if (stb_W_Q0_1_5_0) reg_W_Q0_1_5_0<=wdata[18-1:0];
stb_W_Q0_1_5_1<=(lb.waddr==106)&lb.wren;if (stb_W_Q0_1_5_1) reg_W_Q0_1_5_1<=wdata[18-1:0];
stb_W_Q0_1_5_2<=(lb.waddr==107)&lb.wren;if (stb_W_Q0_1_5_2) reg_W_Q0_1_5_2<=wdata[18-1:0];
stb_W_Q0_1_5_3<=(lb.waddr==108)&lb.wren;if (stb_W_Q0_1_5_3) reg_W_Q0_1_5_3<=wdata[18-1:0];
stb_W_Q0_1_6_0<=(lb.waddr==109)&lb.wren;if (stb_W_Q0_1_6_0) reg_W_Q0_1_6_0<=wdata[18-1:0];
stb_W_Q0_1_6_1<=(lb.waddr==110)&lb.wren;if (stb_W_Q0_1_6_1) reg_W_Q0_1_6_1<=wdata[18-1:0];
stb_W_Q0_1_6_2<=(lb.waddr==111)&lb.wren;if (stb_W_Q0_1_6_2) reg_W_Q0_1_6_2<=wdata[18-1:0];
stb_W_Q0_1_6_3<=(lb.waddr==112)&lb.wren;if (stb_W_Q0_1_6_3) reg_W_Q0_1_6_3<=wdata[18-1:0];
stb_W_Q0_1_7_0<=(lb.waddr==113)&lb.wren;if (stb_W_Q0_1_7_0) reg_W_Q0_1_7_0<=wdata[18-1:0];
stb_W_Q0_1_7_1<=(lb.waddr==114)&lb.wren;if (stb_W_Q0_1_7_1) reg_W_Q0_1_7_1<=wdata[18-1:0];
stb_W_Q0_1_7_2<=(lb.waddr==115)&lb.wren;if (stb_W_Q0_1_7_2) reg_W_Q0_1_7_2<=wdata[18-1:0];
stb_W_Q0_1_7_3<=(lb.waddr==116)&lb.wren;if (stb_W_Q0_1_7_3) reg_W_Q0_1_7_3<=wdata[18-1:0];
stb_W_Q0_2_0_0<=(lb.waddr==117)&lb.wren;if (stb_W_Q0_2_0_0) reg_W_Q0_2_0_0<=wdata[18-1:0];
stb_W_Q0_2_1_0<=(lb.waddr==118)&lb.wren;if (stb_W_Q0_2_1_0) reg_W_Q0_2_1_0<=wdata[18-1:0];
stb_W_Q0_2_2_0<=(lb.waddr==119)&lb.wren;if (stb_W_Q0_2_2_0) reg_W_Q0_2_2_0<=wdata[18-1:0];
stb_W_Q0_2_3_0<=(lb.waddr==120)&lb.wren;if (stb_W_Q0_2_3_0) reg_W_Q0_2_3_0<=wdata[18-1:0];
stb_B_Q0_0_0<=(lb.waddr==121)&lb.wren;if (stb_B_Q0_0_0) reg_B_Q0_0_0<=wdata[18-1:0];
stb_B_Q0_0_1<=(lb.waddr==122)&lb.wren;if (stb_B_Q0_0_1) reg_B_Q0_0_1<=wdata[18-1:0];
stb_B_Q0_0_2<=(lb.waddr==123)&lb.wren;if (stb_B_Q0_0_2) reg_B_Q0_0_2<=wdata[18-1:0];
stb_B_Q0_0_3<=(lb.waddr==124)&lb.wren;if (stb_B_Q0_0_3) reg_B_Q0_0_3<=wdata[18-1:0];
stb_B_Q0_0_4<=(lb.waddr==125)&lb.wren;if (stb_B_Q0_0_4) reg_B_Q0_0_4<=wdata[18-1:0];
stb_B_Q0_0_5<=(lb.waddr==126)&lb.wren;if (stb_B_Q0_0_5) reg_B_Q0_0_5<=wdata[18-1:0];
stb_B_Q0_0_6<=(lb.waddr==127)&lb.wren;if (stb_B_Q0_0_6) reg_B_Q0_0_6<=wdata[18-1:0];
stb_B_Q0_0_7<=(lb.waddr==128)&lb.wren;if (stb_B_Q0_0_7) reg_B_Q0_0_7<=wdata[18-1:0];
stb_B_Q0_1_0<=(lb.waddr==129)&lb.wren;if (stb_B_Q0_1_0) reg_B_Q0_1_0<=wdata[18-1:0];
stb_B_Q0_1_1<=(lb.waddr==130)&lb.wren;if (stb_B_Q0_1_1) reg_B_Q0_1_1<=wdata[18-1:0];
stb_B_Q0_1_2<=(lb.waddr==131)&lb.wren;if (stb_B_Q0_1_2) reg_B_Q0_1_2<=wdata[18-1:0];
stb_B_Q0_1_3<=(lb.waddr==132)&lb.wren;if (stb_B_Q0_1_3) reg_B_Q0_1_3<=wdata[18-1:0];
stb_B_Q0_2_0<=(lb.waddr==133)&lb.wren;if (stb_B_Q0_2_0) reg_B_Q0_2_0<=wdata[18-1:0];
stb_W_Q1_0_0_0<=(lb.waddr==134)&lb.wren;if (stb_W_Q1_0_0_0) reg_W_Q1_0_0_0<=wdata[18-1:0];
stb_W_Q1_0_0_1<=(lb.waddr==135)&lb.wren;if (stb_W_Q1_0_0_1) reg_W_Q1_0_0_1<=wdata[18-1:0];
stb_W_Q1_0_0_2<=(lb.waddr==136)&lb.wren;if (stb_W_Q1_0_0_2) reg_W_Q1_0_0_2<=wdata[18-1:0];
stb_W_Q1_0_0_3<=(lb.waddr==137)&lb.wren;if (stb_W_Q1_0_0_3) reg_W_Q1_0_0_3<=wdata[18-1:0];
stb_W_Q1_0_0_4<=(lb.waddr==138)&lb.wren;if (stb_W_Q1_0_0_4) reg_W_Q1_0_0_4<=wdata[18-1:0];
stb_W_Q1_0_0_5<=(lb.waddr==139)&lb.wren;if (stb_W_Q1_0_0_5) reg_W_Q1_0_0_5<=wdata[18-1:0];
stb_W_Q1_0_0_6<=(lb.waddr==140)&lb.wren;if (stb_W_Q1_0_0_6) reg_W_Q1_0_0_6<=wdata[18-1:0];
stb_W_Q1_0_0_7<=(lb.waddr==141)&lb.wren;if (stb_W_Q1_0_0_7) reg_W_Q1_0_0_7<=wdata[18-1:0];
stb_W_Q1_0_1_0<=(lb.waddr==142)&lb.wren;if (stb_W_Q1_0_1_0) reg_W_Q1_0_1_0<=wdata[18-1:0];
stb_W_Q1_0_1_1<=(lb.waddr==143)&lb.wren;if (stb_W_Q1_0_1_1) reg_W_Q1_0_1_1<=wdata[18-1:0];
stb_W_Q1_0_1_2<=(lb.waddr==144)&lb.wren;if (stb_W_Q1_0_1_2) reg_W_Q1_0_1_2<=wdata[18-1:0];
stb_W_Q1_0_1_3<=(lb.waddr==145)&lb.wren;if (stb_W_Q1_0_1_3) reg_W_Q1_0_1_3<=wdata[18-1:0];
stb_W_Q1_0_1_4<=(lb.waddr==146)&lb.wren;if (stb_W_Q1_0_1_4) reg_W_Q1_0_1_4<=wdata[18-1:0];
stb_W_Q1_0_1_5<=(lb.waddr==147)&lb.wren;if (stb_W_Q1_0_1_5) reg_W_Q1_0_1_5<=wdata[18-1:0];
stb_W_Q1_0_1_6<=(lb.waddr==148)&lb.wren;if (stb_W_Q1_0_1_6) reg_W_Q1_0_1_6<=wdata[18-1:0];
stb_W_Q1_0_1_7<=(lb.waddr==149)&lb.wren;if (stb_W_Q1_0_1_7) reg_W_Q1_0_1_7<=wdata[18-1:0];
stb_W_Q1_1_0_0<=(lb.waddr==150)&lb.wren;if (stb_W_Q1_1_0_0) reg_W_Q1_1_0_0<=wdata[18-1:0];
stb_W_Q1_1_0_1<=(lb.waddr==151)&lb.wren;if (stb_W_Q1_1_0_1) reg_W_Q1_1_0_1<=wdata[18-1:0];
stb_W_Q1_1_0_2<=(lb.waddr==152)&lb.wren;if (stb_W_Q1_1_0_2) reg_W_Q1_1_0_2<=wdata[18-1:0];
stb_W_Q1_1_0_3<=(lb.waddr==153)&lb.wren;if (stb_W_Q1_1_0_3) reg_W_Q1_1_0_3<=wdata[18-1:0];
stb_W_Q1_1_1_0<=(lb.waddr==154)&lb.wren;if (stb_W_Q1_1_1_0) reg_W_Q1_1_1_0<=wdata[18-1:0];
stb_W_Q1_1_1_1<=(lb.waddr==155)&lb.wren;if (stb_W_Q1_1_1_1) reg_W_Q1_1_1_1<=wdata[18-1:0];
stb_W_Q1_1_1_2<=(lb.waddr==156)&lb.wren;if (stb_W_Q1_1_1_2) reg_W_Q1_1_1_2<=wdata[18-1:0];
stb_W_Q1_1_1_3<=(lb.waddr==157)&lb.wren;if (stb_W_Q1_1_1_3) reg_W_Q1_1_1_3<=wdata[18-1:0];
stb_W_Q1_1_2_0<=(lb.waddr==158)&lb.wren;if (stb_W_Q1_1_2_0) reg_W_Q1_1_2_0<=wdata[18-1:0];
stb_W_Q1_1_2_1<=(lb.waddr==159)&lb.wren;if (stb_W_Q1_1_2_1) reg_W_Q1_1_2_1<=wdata[18-1:0];
stb_W_Q1_1_2_2<=(lb.waddr==160)&lb.wren;if (stb_W_Q1_1_2_2) reg_W_Q1_1_2_2<=wdata[18-1:0];
stb_W_Q1_1_2_3<=(lb.waddr==161)&lb.wren;if (stb_W_Q1_1_2_3) reg_W_Q1_1_2_3<=wdata[18-1:0];
stb_W_Q1_1_3_0<=(lb.waddr==162)&lb.wren;if (stb_W_Q1_1_3_0) reg_W_Q1_1_3_0<=wdata[18-1:0];
stb_W_Q1_1_3_1<=(lb.waddr==163)&lb.wren;if (stb_W_Q1_1_3_1) reg_W_Q1_1_3_1<=wdata[18-1:0];
stb_W_Q1_1_3_2<=(lb.waddr==164)&lb.wren;if (stb_W_Q1_1_3_2) reg_W_Q1_1_3_2<=wdata[18-1:0];
stb_W_Q1_1_3_3<=(lb.waddr==165)&lb.wren;if (stb_W_Q1_1_3_3) reg_W_Q1_1_3_3<=wdata[18-1:0];
stb_W_Q1_1_4_0<=(lb.waddr==166)&lb.wren;if (stb_W_Q1_1_4_0) reg_W_Q1_1_4_0<=wdata[18-1:0];
stb_W_Q1_1_4_1<=(lb.waddr==167)&lb.wren;if (stb_W_Q1_1_4_1) reg_W_Q1_1_4_1<=wdata[18-1:0];
stb_W_Q1_1_4_2<=(lb.waddr==168)&lb.wren;if (stb_W_Q1_1_4_2) reg_W_Q1_1_4_2<=wdata[18-1:0];
stb_W_Q1_1_4_3<=(lb.waddr==169)&lb.wren;if (stb_W_Q1_1_4_3) reg_W_Q1_1_4_3<=wdata[18-1:0];
stb_W_Q1_1_5_0<=(lb.waddr==170)&lb.wren;if (stb_W_Q1_1_5_0) reg_W_Q1_1_5_0<=wdata[18-1:0];
stb_W_Q1_1_5_1<=(lb.waddr==171)&lb.wren;if (stb_W_Q1_1_5_1) reg_W_Q1_1_5_1<=wdata[18-1:0];
stb_W_Q1_1_5_2<=(lb.waddr==172)&lb.wren;if (stb_W_Q1_1_5_2) reg_W_Q1_1_5_2<=wdata[18-1:0];
stb_W_Q1_1_5_3<=(lb.waddr==173)&lb.wren;if (stb_W_Q1_1_5_3) reg_W_Q1_1_5_3<=wdata[18-1:0];
stb_W_Q1_1_6_0<=(lb.waddr==174)&lb.wren;if (stb_W_Q1_1_6_0) reg_W_Q1_1_6_0<=wdata[18-1:0];
stb_W_Q1_1_6_1<=(lb.waddr==175)&lb.wren;if (stb_W_Q1_1_6_1) reg_W_Q1_1_6_1<=wdata[18-1:0];
stb_W_Q1_1_6_2<=(lb.waddr==176)&lb.wren;if (stb_W_Q1_1_6_2) reg_W_Q1_1_6_2<=wdata[18-1:0];
stb_W_Q1_1_6_3<=(lb.waddr==177)&lb.wren;if (stb_W_Q1_1_6_3) reg_W_Q1_1_6_3<=wdata[18-1:0];
stb_W_Q1_1_7_0<=(lb.waddr==178)&lb.wren;if (stb_W_Q1_1_7_0) reg_W_Q1_1_7_0<=wdata[18-1:0];
stb_W_Q1_1_7_1<=(lb.waddr==179)&lb.wren;if (stb_W_Q1_1_7_1) reg_W_Q1_1_7_1<=wdata[18-1:0];
stb_W_Q1_1_7_2<=(lb.waddr==180)&lb.wren;if (stb_W_Q1_1_7_2) reg_W_Q1_1_7_2<=wdata[18-1:0];
stb_W_Q1_1_7_3<=(lb.waddr==181)&lb.wren;if (stb_W_Q1_1_7_3) reg_W_Q1_1_7_3<=wdata[18-1:0];
stb_W_Q1_2_0_0<=(lb.waddr==182)&lb.wren;if (stb_W_Q1_2_0_0) reg_W_Q1_2_0_0<=wdata[18-1:0];
stb_W_Q1_2_1_0<=(lb.waddr==183)&lb.wren;if (stb_W_Q1_2_1_0) reg_W_Q1_2_1_0<=wdata[18-1:0];
stb_W_Q1_2_2_0<=(lb.waddr==184)&lb.wren;if (stb_W_Q1_2_2_0) reg_W_Q1_2_2_0<=wdata[18-1:0];
stb_W_Q1_2_3_0<=(lb.waddr==185)&lb.wren;if (stb_W_Q1_2_3_0) reg_W_Q1_2_3_0<=wdata[18-1:0];
stb_B_Q1_0_0<=(lb.waddr==186)&lb.wren;if (stb_B_Q1_0_0) reg_B_Q1_0_0<=wdata[18-1:0];
stb_B_Q1_0_1<=(lb.waddr==187)&lb.wren;if (stb_B_Q1_0_1) reg_B_Q1_0_1<=wdata[18-1:0];
stb_B_Q1_0_2<=(lb.waddr==188)&lb.wren;if (stb_B_Q1_0_2) reg_B_Q1_0_2<=wdata[18-1:0];
stb_B_Q1_0_3<=(lb.waddr==189)&lb.wren;if (stb_B_Q1_0_3) reg_B_Q1_0_3<=wdata[18-1:0];
stb_B_Q1_0_4<=(lb.waddr==190)&lb.wren;if (stb_B_Q1_0_4) reg_B_Q1_0_4<=wdata[18-1:0];
stb_B_Q1_0_5<=(lb.waddr==191)&lb.wren;if (stb_B_Q1_0_5) reg_B_Q1_0_5<=wdata[18-1:0];
stb_B_Q1_0_6<=(lb.waddr==192)&lb.wren;if (stb_B_Q1_0_6) reg_B_Q1_0_6<=wdata[18-1:0];
stb_B_Q1_0_7<=(lb.waddr==193)&lb.wren;if (stb_B_Q1_0_7) reg_B_Q1_0_7<=wdata[18-1:0];
stb_B_Q1_1_0<=(lb.waddr==194)&lb.wren;if (stb_B_Q1_1_0) reg_B_Q1_1_0<=wdata[18-1:0];
stb_B_Q1_1_1<=(lb.waddr==195)&lb.wren;if (stb_B_Q1_1_1) reg_B_Q1_1_1<=wdata[18-1:0];
stb_B_Q1_1_2<=(lb.waddr==196)&lb.wren;if (stb_B_Q1_1_2) reg_B_Q1_1_2<=wdata[18-1:0];
stb_B_Q1_1_3<=(lb.waddr==197)&lb.wren;if (stb_B_Q1_1_3) reg_B_Q1_1_3<=wdata[18-1:0];
stb_B_Q1_2_0<=(lb.waddr==198)&lb.wren;if (stb_B_Q1_2_0) reg_B_Q1_2_0<=wdata[18-1:0];
stb_W_Q2_0_0_0<=(lb.waddr==199)&lb.wren;if (stb_W_Q2_0_0_0) reg_W_Q2_0_0_0<=wdata[18-1:0];
stb_W_Q2_0_0_1<=(lb.waddr==200)&lb.wren;if (stb_W_Q2_0_0_1) reg_W_Q2_0_0_1<=wdata[18-1:0];
stb_W_Q2_0_0_2<=(lb.waddr==201)&lb.wren;if (stb_W_Q2_0_0_2) reg_W_Q2_0_0_2<=wdata[18-1:0];
stb_W_Q2_0_0_3<=(lb.waddr==202)&lb.wren;if (stb_W_Q2_0_0_3) reg_W_Q2_0_0_3<=wdata[18-1:0];
stb_W_Q2_0_0_4<=(lb.waddr==203)&lb.wren;if (stb_W_Q2_0_0_4) reg_W_Q2_0_0_4<=wdata[18-1:0];
stb_W_Q2_0_0_5<=(lb.waddr==204)&lb.wren;if (stb_W_Q2_0_0_5) reg_W_Q2_0_0_5<=wdata[18-1:0];
stb_W_Q2_0_0_6<=(lb.waddr==205)&lb.wren;if (stb_W_Q2_0_0_6) reg_W_Q2_0_0_6<=wdata[18-1:0];
stb_W_Q2_0_0_7<=(lb.waddr==206)&lb.wren;if (stb_W_Q2_0_0_7) reg_W_Q2_0_0_7<=wdata[18-1:0];
stb_W_Q2_0_1_0<=(lb.waddr==207)&lb.wren;if (stb_W_Q2_0_1_0) reg_W_Q2_0_1_0<=wdata[18-1:0];
stb_W_Q2_0_1_1<=(lb.waddr==208)&lb.wren;if (stb_W_Q2_0_1_1) reg_W_Q2_0_1_1<=wdata[18-1:0];
stb_W_Q2_0_1_2<=(lb.waddr==209)&lb.wren;if (stb_W_Q2_0_1_2) reg_W_Q2_0_1_2<=wdata[18-1:0];
stb_W_Q2_0_1_3<=(lb.waddr==210)&lb.wren;if (stb_W_Q2_0_1_3) reg_W_Q2_0_1_3<=wdata[18-1:0];
stb_W_Q2_0_1_4<=(lb.waddr==211)&lb.wren;if (stb_W_Q2_0_1_4) reg_W_Q2_0_1_4<=wdata[18-1:0];
stb_W_Q2_0_1_5<=(lb.waddr==212)&lb.wren;if (stb_W_Q2_0_1_5) reg_W_Q2_0_1_5<=wdata[18-1:0];
stb_W_Q2_0_1_6<=(lb.waddr==213)&lb.wren;if (stb_W_Q2_0_1_6) reg_W_Q2_0_1_6<=wdata[18-1:0];
stb_W_Q2_0_1_7<=(lb.waddr==214)&lb.wren;if (stb_W_Q2_0_1_7) reg_W_Q2_0_1_7<=wdata[18-1:0];
stb_W_Q2_1_0_0<=(lb.waddr==215)&lb.wren;if (stb_W_Q2_1_0_0) reg_W_Q2_1_0_0<=wdata[18-1:0];
stb_W_Q2_1_0_1<=(lb.waddr==216)&lb.wren;if (stb_W_Q2_1_0_1) reg_W_Q2_1_0_1<=wdata[18-1:0];
stb_W_Q2_1_0_2<=(lb.waddr==217)&lb.wren;if (stb_W_Q2_1_0_2) reg_W_Q2_1_0_2<=wdata[18-1:0];
stb_W_Q2_1_0_3<=(lb.waddr==218)&lb.wren;if (stb_W_Q2_1_0_3) reg_W_Q2_1_0_3<=wdata[18-1:0];
stb_W_Q2_1_1_0<=(lb.waddr==219)&lb.wren;if (stb_W_Q2_1_1_0) reg_W_Q2_1_1_0<=wdata[18-1:0];
stb_W_Q2_1_1_1<=(lb.waddr==220)&lb.wren;if (stb_W_Q2_1_1_1) reg_W_Q2_1_1_1<=wdata[18-1:0];
stb_W_Q2_1_1_2<=(lb.waddr==221)&lb.wren;if (stb_W_Q2_1_1_2) reg_W_Q2_1_1_2<=wdata[18-1:0];
stb_W_Q2_1_1_3<=(lb.waddr==222)&lb.wren;if (stb_W_Q2_1_1_3) reg_W_Q2_1_1_3<=wdata[18-1:0];
stb_W_Q2_1_2_0<=(lb.waddr==223)&lb.wren;if (stb_W_Q2_1_2_0) reg_W_Q2_1_2_0<=wdata[18-1:0];
stb_W_Q2_1_2_1<=(lb.waddr==224)&lb.wren;if (stb_W_Q2_1_2_1) reg_W_Q2_1_2_1<=wdata[18-1:0];
stb_W_Q2_1_2_2<=(lb.waddr==225)&lb.wren;if (stb_W_Q2_1_2_2) reg_W_Q2_1_2_2<=wdata[18-1:0];
stb_W_Q2_1_2_3<=(lb.waddr==226)&lb.wren;if (stb_W_Q2_1_2_3) reg_W_Q2_1_2_3<=wdata[18-1:0];
stb_W_Q2_1_3_0<=(lb.waddr==227)&lb.wren;if (stb_W_Q2_1_3_0) reg_W_Q2_1_3_0<=wdata[18-1:0];
stb_W_Q2_1_3_1<=(lb.waddr==228)&lb.wren;if (stb_W_Q2_1_3_1) reg_W_Q2_1_3_1<=wdata[18-1:0];
stb_W_Q2_1_3_2<=(lb.waddr==229)&lb.wren;if (stb_W_Q2_1_3_2) reg_W_Q2_1_3_2<=wdata[18-1:0];
stb_W_Q2_1_3_3<=(lb.waddr==230)&lb.wren;if (stb_W_Q2_1_3_3) reg_W_Q2_1_3_3<=wdata[18-1:0];
stb_W_Q2_1_4_0<=(lb.waddr==231)&lb.wren;if (stb_W_Q2_1_4_0) reg_W_Q2_1_4_0<=wdata[18-1:0];
stb_W_Q2_1_4_1<=(lb.waddr==232)&lb.wren;if (stb_W_Q2_1_4_1) reg_W_Q2_1_4_1<=wdata[18-1:0];
stb_W_Q2_1_4_2<=(lb.waddr==233)&lb.wren;if (stb_W_Q2_1_4_2) reg_W_Q2_1_4_2<=wdata[18-1:0];
stb_W_Q2_1_4_3<=(lb.waddr==234)&lb.wren;if (stb_W_Q2_1_4_3) reg_W_Q2_1_4_3<=wdata[18-1:0];
stb_W_Q2_1_5_0<=(lb.waddr==235)&lb.wren;if (stb_W_Q2_1_5_0) reg_W_Q2_1_5_0<=wdata[18-1:0];
stb_W_Q2_1_5_1<=(lb.waddr==236)&lb.wren;if (stb_W_Q2_1_5_1) reg_W_Q2_1_5_1<=wdata[18-1:0];
stb_W_Q2_1_5_2<=(lb.waddr==237)&lb.wren;if (stb_W_Q2_1_5_2) reg_W_Q2_1_5_2<=wdata[18-1:0];
stb_W_Q2_1_5_3<=(lb.waddr==238)&lb.wren;if (stb_W_Q2_1_5_3) reg_W_Q2_1_5_3<=wdata[18-1:0];
stb_W_Q2_1_6_0<=(lb.waddr==239)&lb.wren;if (stb_W_Q2_1_6_0) reg_W_Q2_1_6_0<=wdata[18-1:0];
stb_W_Q2_1_6_1<=(lb.waddr==240)&lb.wren;if (stb_W_Q2_1_6_1) reg_W_Q2_1_6_1<=wdata[18-1:0];
stb_W_Q2_1_6_2<=(lb.waddr==241)&lb.wren;if (stb_W_Q2_1_6_2) reg_W_Q2_1_6_2<=wdata[18-1:0];
stb_W_Q2_1_6_3<=(lb.waddr==242)&lb.wren;if (stb_W_Q2_1_6_3) reg_W_Q2_1_6_3<=wdata[18-1:0];
stb_W_Q2_1_7_0<=(lb.waddr==243)&lb.wren;if (stb_W_Q2_1_7_0) reg_W_Q2_1_7_0<=wdata[18-1:0];
stb_W_Q2_1_7_1<=(lb.waddr==244)&lb.wren;if (stb_W_Q2_1_7_1) reg_W_Q2_1_7_1<=wdata[18-1:0];
stb_W_Q2_1_7_2<=(lb.waddr==245)&lb.wren;if (stb_W_Q2_1_7_2) reg_W_Q2_1_7_2<=wdata[18-1:0];
stb_W_Q2_1_7_3<=(lb.waddr==246)&lb.wren;if (stb_W_Q2_1_7_3) reg_W_Q2_1_7_3<=wdata[18-1:0];
stb_W_Q2_2_0_0<=(lb.waddr==247)&lb.wren;if (stb_W_Q2_2_0_0) reg_W_Q2_2_0_0<=wdata[18-1:0];
stb_W_Q2_2_1_0<=(lb.waddr==248)&lb.wren;if (stb_W_Q2_2_1_0) reg_W_Q2_2_1_0<=wdata[18-1:0];
stb_W_Q2_2_2_0<=(lb.waddr==249)&lb.wren;if (stb_W_Q2_2_2_0) reg_W_Q2_2_2_0<=wdata[18-1:0];
stb_W_Q2_2_3_0<=(lb.waddr==250)&lb.wren;if (stb_W_Q2_2_3_0) reg_W_Q2_2_3_0<=wdata[18-1:0];
stb_B_Q2_0_0<=(lb.waddr==251)&lb.wren;if (stb_B_Q2_0_0) reg_B_Q2_0_0<=wdata[18-1:0];
stb_B_Q2_0_1<=(lb.waddr==252)&lb.wren;if (stb_B_Q2_0_1) reg_B_Q2_0_1<=wdata[18-1:0];
stb_B_Q2_0_2<=(lb.waddr==253)&lb.wren;if (stb_B_Q2_0_2) reg_B_Q2_0_2<=wdata[18-1:0];
stb_B_Q2_0_3<=(lb.waddr==254)&lb.wren;if (stb_B_Q2_0_3) reg_B_Q2_0_3<=wdata[18-1:0];
stb_B_Q2_0_4<=(lb.waddr==255)&lb.wren;if (stb_B_Q2_0_4) reg_B_Q2_0_4<=wdata[18-1:0];
stb_B_Q2_0_5<=(lb.waddr==256)&lb.wren;if (stb_B_Q2_0_5) reg_B_Q2_0_5<=wdata[18-1:0];
stb_B_Q2_0_6<=(lb.waddr==257)&lb.wren;if (stb_B_Q2_0_6) reg_B_Q2_0_6<=wdata[18-1:0];
stb_B_Q2_0_7<=(lb.waddr==258)&lb.wren;if (stb_B_Q2_0_7) reg_B_Q2_0_7<=wdata[18-1:0];
stb_B_Q2_1_0<=(lb.waddr==259)&lb.wren;if (stb_B_Q2_1_0) reg_B_Q2_1_0<=wdata[18-1:0];
stb_B_Q2_1_1<=(lb.waddr==260)&lb.wren;if (stb_B_Q2_1_1) reg_B_Q2_1_1<=wdata[18-1:0];
stb_B_Q2_1_2<=(lb.waddr==261)&lb.wren;if (stb_B_Q2_1_2) reg_B_Q2_1_2<=wdata[18-1:0];
stb_B_Q2_1_3<=(lb.waddr==262)&lb.wren;if (stb_B_Q2_1_3) reg_B_Q2_1_3<=wdata[18-1:0];
stb_B_Q2_2_0<=(lb.waddr==263)&lb.wren;if (stb_B_Q2_2_0) reg_B_Q2_2_0<=wdata[18-1:0];
stb_W_Q3_0_0_0<=(lb.waddr==264)&lb.wren;if (stb_W_Q3_0_0_0) reg_W_Q3_0_0_0<=wdata[18-1:0];
stb_W_Q3_0_0_1<=(lb.waddr==265)&lb.wren;if (stb_W_Q3_0_0_1) reg_W_Q3_0_0_1<=wdata[18-1:0];
stb_W_Q3_0_0_2<=(lb.waddr==266)&lb.wren;if (stb_W_Q3_0_0_2) reg_W_Q3_0_0_2<=wdata[18-1:0];
stb_W_Q3_0_0_3<=(lb.waddr==267)&lb.wren;if (stb_W_Q3_0_0_3) reg_W_Q3_0_0_3<=wdata[18-1:0];
stb_W_Q3_0_0_4<=(lb.waddr==268)&lb.wren;if (stb_W_Q3_0_0_4) reg_W_Q3_0_0_4<=wdata[18-1:0];
stb_W_Q3_0_0_5<=(lb.waddr==269)&lb.wren;if (stb_W_Q3_0_0_5) reg_W_Q3_0_0_5<=wdata[18-1:0];
stb_W_Q3_0_0_6<=(lb.waddr==270)&lb.wren;if (stb_W_Q3_0_0_6) reg_W_Q3_0_0_6<=wdata[18-1:0];
stb_W_Q3_0_0_7<=(lb.waddr==271)&lb.wren;if (stb_W_Q3_0_0_7) reg_W_Q3_0_0_7<=wdata[18-1:0];
stb_W_Q3_0_1_0<=(lb.waddr==272)&lb.wren;if (stb_W_Q3_0_1_0) reg_W_Q3_0_1_0<=wdata[18-1:0];
stb_W_Q3_0_1_1<=(lb.waddr==273)&lb.wren;if (stb_W_Q3_0_1_1) reg_W_Q3_0_1_1<=wdata[18-1:0];
stb_W_Q3_0_1_2<=(lb.waddr==274)&lb.wren;if (stb_W_Q3_0_1_2) reg_W_Q3_0_1_2<=wdata[18-1:0];
stb_W_Q3_0_1_3<=(lb.waddr==275)&lb.wren;if (stb_W_Q3_0_1_3) reg_W_Q3_0_1_3<=wdata[18-1:0];
stb_W_Q3_0_1_4<=(lb.waddr==276)&lb.wren;if (stb_W_Q3_0_1_4) reg_W_Q3_0_1_4<=wdata[18-1:0];
stb_W_Q3_0_1_5<=(lb.waddr==277)&lb.wren;if (stb_W_Q3_0_1_5) reg_W_Q3_0_1_5<=wdata[18-1:0];
stb_W_Q3_0_1_6<=(lb.waddr==278)&lb.wren;if (stb_W_Q3_0_1_6) reg_W_Q3_0_1_6<=wdata[18-1:0];
stb_W_Q3_0_1_7<=(lb.waddr==279)&lb.wren;if (stb_W_Q3_0_1_7) reg_W_Q3_0_1_7<=wdata[18-1:0];
stb_W_Q3_1_0_0<=(lb.waddr==280)&lb.wren;if (stb_W_Q3_1_0_0) reg_W_Q3_1_0_0<=wdata[18-1:0];
stb_W_Q3_1_0_1<=(lb.waddr==281)&lb.wren;if (stb_W_Q3_1_0_1) reg_W_Q3_1_0_1<=wdata[18-1:0];
stb_W_Q3_1_0_2<=(lb.waddr==282)&lb.wren;if (stb_W_Q3_1_0_2) reg_W_Q3_1_0_2<=wdata[18-1:0];
stb_W_Q3_1_0_3<=(lb.waddr==283)&lb.wren;if (stb_W_Q3_1_0_3) reg_W_Q3_1_0_3<=wdata[18-1:0];
stb_W_Q3_1_1_0<=(lb.waddr==284)&lb.wren;if (stb_W_Q3_1_1_0) reg_W_Q3_1_1_0<=wdata[18-1:0];
stb_W_Q3_1_1_1<=(lb.waddr==285)&lb.wren;if (stb_W_Q3_1_1_1) reg_W_Q3_1_1_1<=wdata[18-1:0];
stb_W_Q3_1_1_2<=(lb.waddr==286)&lb.wren;if (stb_W_Q3_1_1_2) reg_W_Q3_1_1_2<=wdata[18-1:0];
stb_W_Q3_1_1_3<=(lb.waddr==287)&lb.wren;if (stb_W_Q3_1_1_3) reg_W_Q3_1_1_3<=wdata[18-1:0];
stb_W_Q3_1_2_0<=(lb.waddr==288)&lb.wren;if (stb_W_Q3_1_2_0) reg_W_Q3_1_2_0<=wdata[18-1:0];
stb_W_Q3_1_2_1<=(lb.waddr==289)&lb.wren;if (stb_W_Q3_1_2_1) reg_W_Q3_1_2_1<=wdata[18-1:0];
stb_W_Q3_1_2_2<=(lb.waddr==290)&lb.wren;if (stb_W_Q3_1_2_2) reg_W_Q3_1_2_2<=wdata[18-1:0];
stb_W_Q3_1_2_3<=(lb.waddr==291)&lb.wren;if (stb_W_Q3_1_2_3) reg_W_Q3_1_2_3<=wdata[18-1:0];
stb_W_Q3_1_3_0<=(lb.waddr==292)&lb.wren;if (stb_W_Q3_1_3_0) reg_W_Q3_1_3_0<=wdata[18-1:0];
stb_W_Q3_1_3_1<=(lb.waddr==293)&lb.wren;if (stb_W_Q3_1_3_1) reg_W_Q3_1_3_1<=wdata[18-1:0];
stb_W_Q3_1_3_2<=(lb.waddr==294)&lb.wren;if (stb_W_Q3_1_3_2) reg_W_Q3_1_3_2<=wdata[18-1:0];
stb_W_Q3_1_3_3<=(lb.waddr==295)&lb.wren;if (stb_W_Q3_1_3_3) reg_W_Q3_1_3_3<=wdata[18-1:0];
stb_W_Q3_1_4_0<=(lb.waddr==296)&lb.wren;if (stb_W_Q3_1_4_0) reg_W_Q3_1_4_0<=wdata[18-1:0];
stb_W_Q3_1_4_1<=(lb.waddr==297)&lb.wren;if (stb_W_Q3_1_4_1) reg_W_Q3_1_4_1<=wdata[18-1:0];
stb_W_Q3_1_4_2<=(lb.waddr==298)&lb.wren;if (stb_W_Q3_1_4_2) reg_W_Q3_1_4_2<=wdata[18-1:0];
stb_W_Q3_1_4_3<=(lb.waddr==299)&lb.wren;if (stb_W_Q3_1_4_3) reg_W_Q3_1_4_3<=wdata[18-1:0];
stb_W_Q3_1_5_0<=(lb.waddr==300)&lb.wren;if (stb_W_Q3_1_5_0) reg_W_Q3_1_5_0<=wdata[18-1:0];
stb_W_Q3_1_5_1<=(lb.waddr==301)&lb.wren;if (stb_W_Q3_1_5_1) reg_W_Q3_1_5_1<=wdata[18-1:0];
stb_W_Q3_1_5_2<=(lb.waddr==302)&lb.wren;if (stb_W_Q3_1_5_2) reg_W_Q3_1_5_2<=wdata[18-1:0];
stb_W_Q3_1_5_3<=(lb.waddr==303)&lb.wren;if (stb_W_Q3_1_5_3) reg_W_Q3_1_5_3<=wdata[18-1:0];
stb_W_Q3_1_6_0<=(lb.waddr==304)&lb.wren;if (stb_W_Q3_1_6_0) reg_W_Q3_1_6_0<=wdata[18-1:0];
stb_W_Q3_1_6_1<=(lb.waddr==305)&lb.wren;if (stb_W_Q3_1_6_1) reg_W_Q3_1_6_1<=wdata[18-1:0];
stb_W_Q3_1_6_2<=(lb.waddr==306)&lb.wren;if (stb_W_Q3_1_6_2) reg_W_Q3_1_6_2<=wdata[18-1:0];
stb_W_Q3_1_6_3<=(lb.waddr==307)&lb.wren;if (stb_W_Q3_1_6_3) reg_W_Q3_1_6_3<=wdata[18-1:0];
stb_W_Q3_1_7_0<=(lb.waddr==308)&lb.wren;if (stb_W_Q3_1_7_0) reg_W_Q3_1_7_0<=wdata[18-1:0];
stb_W_Q3_1_7_1<=(lb.waddr==309)&lb.wren;if (stb_W_Q3_1_7_1) reg_W_Q3_1_7_1<=wdata[18-1:0];
stb_W_Q3_1_7_2<=(lb.waddr==310)&lb.wren;if (stb_W_Q3_1_7_2) reg_W_Q3_1_7_2<=wdata[18-1:0];
stb_W_Q3_1_7_3<=(lb.waddr==311)&lb.wren;if (stb_W_Q3_1_7_3) reg_W_Q3_1_7_3<=wdata[18-1:0];
stb_W_Q3_2_0_0<=(lb.waddr==312)&lb.wren;if (stb_W_Q3_2_0_0) reg_W_Q3_2_0_0<=wdata[18-1:0];
stb_W_Q3_2_1_0<=(lb.waddr==313)&lb.wren;if (stb_W_Q3_2_1_0) reg_W_Q3_2_1_0<=wdata[18-1:0];
stb_W_Q3_2_2_0<=(lb.waddr==314)&lb.wren;if (stb_W_Q3_2_2_0) reg_W_Q3_2_2_0<=wdata[18-1:0];
stb_W_Q3_2_3_0<=(lb.waddr==315)&lb.wren;if (stb_W_Q3_2_3_0) reg_W_Q3_2_3_0<=wdata[18-1:0];
stb_B_Q3_0_0<=(lb.waddr==316)&lb.wren;if (stb_B_Q3_0_0) reg_B_Q3_0_0<=wdata[18-1:0];
stb_B_Q3_0_1<=(lb.waddr==317)&lb.wren;if (stb_B_Q3_0_1) reg_B_Q3_0_1<=wdata[18-1:0];
stb_B_Q3_0_2<=(lb.waddr==318)&lb.wren;if (stb_B_Q3_0_2) reg_B_Q3_0_2<=wdata[18-1:0];
stb_B_Q3_0_3<=(lb.waddr==319)&lb.wren;if (stb_B_Q3_0_3) reg_B_Q3_0_3<=wdata[18-1:0];
stb_B_Q3_0_4<=(lb.waddr==320)&lb.wren;if (stb_B_Q3_0_4) reg_B_Q3_0_4<=wdata[18-1:0];
stb_B_Q3_0_5<=(lb.waddr==321)&lb.wren;if (stb_B_Q3_0_5) reg_B_Q3_0_5<=wdata[18-1:0];
stb_B_Q3_0_6<=(lb.waddr==322)&lb.wren;if (stb_B_Q3_0_6) reg_B_Q3_0_6<=wdata[18-1:0];
stb_B_Q3_0_7<=(lb.waddr==323)&lb.wren;if (stb_B_Q3_0_7) reg_B_Q3_0_7<=wdata[18-1:0];
stb_B_Q3_1_0<=(lb.waddr==324)&lb.wren;if (stb_B_Q3_1_0) reg_B_Q3_1_0<=wdata[18-1:0];
stb_B_Q3_1_1<=(lb.waddr==325)&lb.wren;if (stb_B_Q3_1_1) reg_B_Q3_1_1<=wdata[18-1:0];
stb_B_Q3_1_2<=(lb.waddr==326)&lb.wren;if (stb_B_Q3_1_2) reg_B_Q3_1_2<=wdata[18-1:0];
stb_B_Q3_1_3<=(lb.waddr==327)&lb.wren;if (stb_B_Q3_1_3) reg_B_Q3_1_3<=wdata[18-1:0];
stb_B_Q3_2_0<=(lb.waddr==328)&lb.wren;if (stb_B_Q3_2_0) reg_B_Q3_2_0<=wdata[18-1:0];
stb_W_Q4_0_0_0<=(lb.waddr==329)&lb.wren;if (stb_W_Q4_0_0_0) reg_W_Q4_0_0_0<=wdata[18-1:0];
stb_W_Q4_0_0_1<=(lb.waddr==330)&lb.wren;if (stb_W_Q4_0_0_1) reg_W_Q4_0_0_1<=wdata[18-1:0];
stb_W_Q4_0_0_2<=(lb.waddr==331)&lb.wren;if (stb_W_Q4_0_0_2) reg_W_Q4_0_0_2<=wdata[18-1:0];
stb_W_Q4_0_0_3<=(lb.waddr==332)&lb.wren;if (stb_W_Q4_0_0_3) reg_W_Q4_0_0_3<=wdata[18-1:0];
stb_W_Q4_0_0_4<=(lb.waddr==333)&lb.wren;if (stb_W_Q4_0_0_4) reg_W_Q4_0_0_4<=wdata[18-1:0];
stb_W_Q4_0_0_5<=(lb.waddr==334)&lb.wren;if (stb_W_Q4_0_0_5) reg_W_Q4_0_0_5<=wdata[18-1:0];
stb_W_Q4_0_0_6<=(lb.waddr==335)&lb.wren;if (stb_W_Q4_0_0_6) reg_W_Q4_0_0_6<=wdata[18-1:0];
stb_W_Q4_0_0_7<=(lb.waddr==336)&lb.wren;if (stb_W_Q4_0_0_7) reg_W_Q4_0_0_7<=wdata[18-1:0];
stb_W_Q4_0_1_0<=(lb.waddr==337)&lb.wren;if (stb_W_Q4_0_1_0) reg_W_Q4_0_1_0<=wdata[18-1:0];
stb_W_Q4_0_1_1<=(lb.waddr==338)&lb.wren;if (stb_W_Q4_0_1_1) reg_W_Q4_0_1_1<=wdata[18-1:0];
stb_W_Q4_0_1_2<=(lb.waddr==339)&lb.wren;if (stb_W_Q4_0_1_2) reg_W_Q4_0_1_2<=wdata[18-1:0];
stb_W_Q4_0_1_3<=(lb.waddr==340)&lb.wren;if (stb_W_Q4_0_1_3) reg_W_Q4_0_1_3<=wdata[18-1:0];
stb_W_Q4_0_1_4<=(lb.waddr==341)&lb.wren;if (stb_W_Q4_0_1_4) reg_W_Q4_0_1_4<=wdata[18-1:0];
stb_W_Q4_0_1_5<=(lb.waddr==342)&lb.wren;if (stb_W_Q4_0_1_5) reg_W_Q4_0_1_5<=wdata[18-1:0];
stb_W_Q4_0_1_6<=(lb.waddr==343)&lb.wren;if (stb_W_Q4_0_1_6) reg_W_Q4_0_1_6<=wdata[18-1:0];
stb_W_Q4_0_1_7<=(lb.waddr==344)&lb.wren;if (stb_W_Q4_0_1_7) reg_W_Q4_0_1_7<=wdata[18-1:0];
stb_W_Q4_1_0_0<=(lb.waddr==345)&lb.wren;if (stb_W_Q4_1_0_0) reg_W_Q4_1_0_0<=wdata[18-1:0];
stb_W_Q4_1_0_1<=(lb.waddr==346)&lb.wren;if (stb_W_Q4_1_0_1) reg_W_Q4_1_0_1<=wdata[18-1:0];
stb_W_Q4_1_0_2<=(lb.waddr==347)&lb.wren;if (stb_W_Q4_1_0_2) reg_W_Q4_1_0_2<=wdata[18-1:0];
stb_W_Q4_1_0_3<=(lb.waddr==348)&lb.wren;if (stb_W_Q4_1_0_3) reg_W_Q4_1_0_3<=wdata[18-1:0];
stb_W_Q4_1_1_0<=(lb.waddr==349)&lb.wren;if (stb_W_Q4_1_1_0) reg_W_Q4_1_1_0<=wdata[18-1:0];
stb_W_Q4_1_1_1<=(lb.waddr==350)&lb.wren;if (stb_W_Q4_1_1_1) reg_W_Q4_1_1_1<=wdata[18-1:0];
stb_W_Q4_1_1_2<=(lb.waddr==351)&lb.wren;if (stb_W_Q4_1_1_2) reg_W_Q4_1_1_2<=wdata[18-1:0];
stb_W_Q4_1_1_3<=(lb.waddr==352)&lb.wren;if (stb_W_Q4_1_1_3) reg_W_Q4_1_1_3<=wdata[18-1:0];
stb_W_Q4_1_2_0<=(lb.waddr==353)&lb.wren;if (stb_W_Q4_1_2_0) reg_W_Q4_1_2_0<=wdata[18-1:0];
stb_W_Q4_1_2_1<=(lb.waddr==354)&lb.wren;if (stb_W_Q4_1_2_1) reg_W_Q4_1_2_1<=wdata[18-1:0];
stb_W_Q4_1_2_2<=(lb.waddr==355)&lb.wren;if (stb_W_Q4_1_2_2) reg_W_Q4_1_2_2<=wdata[18-1:0];
stb_W_Q4_1_2_3<=(lb.waddr==356)&lb.wren;if (stb_W_Q4_1_2_3) reg_W_Q4_1_2_3<=wdata[18-1:0];
stb_W_Q4_1_3_0<=(lb.waddr==357)&lb.wren;if (stb_W_Q4_1_3_0) reg_W_Q4_1_3_0<=wdata[18-1:0];
stb_W_Q4_1_3_1<=(lb.waddr==358)&lb.wren;if (stb_W_Q4_1_3_1) reg_W_Q4_1_3_1<=wdata[18-1:0];
stb_W_Q4_1_3_2<=(lb.waddr==359)&lb.wren;if (stb_W_Q4_1_3_2) reg_W_Q4_1_3_2<=wdata[18-1:0];
stb_W_Q4_1_3_3<=(lb.waddr==360)&lb.wren;if (stb_W_Q4_1_3_3) reg_W_Q4_1_3_3<=wdata[18-1:0];
stb_W_Q4_1_4_0<=(lb.waddr==361)&lb.wren;if (stb_W_Q4_1_4_0) reg_W_Q4_1_4_0<=wdata[18-1:0];
stb_W_Q4_1_4_1<=(lb.waddr==362)&lb.wren;if (stb_W_Q4_1_4_1) reg_W_Q4_1_4_1<=wdata[18-1:0];
stb_W_Q4_1_4_2<=(lb.waddr==363)&lb.wren;if (stb_W_Q4_1_4_2) reg_W_Q4_1_4_2<=wdata[18-1:0];
stb_W_Q4_1_4_3<=(lb.waddr==364)&lb.wren;if (stb_W_Q4_1_4_3) reg_W_Q4_1_4_3<=wdata[18-1:0];
stb_W_Q4_1_5_0<=(lb.waddr==365)&lb.wren;if (stb_W_Q4_1_5_0) reg_W_Q4_1_5_0<=wdata[18-1:0];
stb_W_Q4_1_5_1<=(lb.waddr==366)&lb.wren;if (stb_W_Q4_1_5_1) reg_W_Q4_1_5_1<=wdata[18-1:0];
stb_W_Q4_1_5_2<=(lb.waddr==367)&lb.wren;if (stb_W_Q4_1_5_2) reg_W_Q4_1_5_2<=wdata[18-1:0];
stb_W_Q4_1_5_3<=(lb.waddr==368)&lb.wren;if (stb_W_Q4_1_5_3) reg_W_Q4_1_5_3<=wdata[18-1:0];
stb_W_Q4_1_6_0<=(lb.waddr==369)&lb.wren;if (stb_W_Q4_1_6_0) reg_W_Q4_1_6_0<=wdata[18-1:0];
stb_W_Q4_1_6_1<=(lb.waddr==370)&lb.wren;if (stb_W_Q4_1_6_1) reg_W_Q4_1_6_1<=wdata[18-1:0];
stb_W_Q4_1_6_2<=(lb.waddr==371)&lb.wren;if (stb_W_Q4_1_6_2) reg_W_Q4_1_6_2<=wdata[18-1:0];
stb_W_Q4_1_6_3<=(lb.waddr==372)&lb.wren;if (stb_W_Q4_1_6_3) reg_W_Q4_1_6_3<=wdata[18-1:0];
stb_W_Q4_1_7_0<=(lb.waddr==373)&lb.wren;if (stb_W_Q4_1_7_0) reg_W_Q4_1_7_0<=wdata[18-1:0];
stb_W_Q4_1_7_1<=(lb.waddr==374)&lb.wren;if (stb_W_Q4_1_7_1) reg_W_Q4_1_7_1<=wdata[18-1:0];
stb_W_Q4_1_7_2<=(lb.waddr==375)&lb.wren;if (stb_W_Q4_1_7_2) reg_W_Q4_1_7_2<=wdata[18-1:0];
stb_W_Q4_1_7_3<=(lb.waddr==376)&lb.wren;if (stb_W_Q4_1_7_3) reg_W_Q4_1_7_3<=wdata[18-1:0];
stb_W_Q4_2_0_0<=(lb.waddr==377)&lb.wren;if (stb_W_Q4_2_0_0) reg_W_Q4_2_0_0<=wdata[18-1:0];
stb_W_Q4_2_1_0<=(lb.waddr==378)&lb.wren;if (stb_W_Q4_2_1_0) reg_W_Q4_2_1_0<=wdata[18-1:0];
stb_W_Q4_2_2_0<=(lb.waddr==379)&lb.wren;if (stb_W_Q4_2_2_0) reg_W_Q4_2_2_0<=wdata[18-1:0];
stb_W_Q4_2_3_0<=(lb.waddr==380)&lb.wren;if (stb_W_Q4_2_3_0) reg_W_Q4_2_3_0<=wdata[18-1:0];
stb_B_Q4_0_0<=(lb.waddr==381)&lb.wren;if (stb_B_Q4_0_0) reg_B_Q4_0_0<=wdata[18-1:0];
stb_B_Q4_0_1<=(lb.waddr==382)&lb.wren;if (stb_B_Q4_0_1) reg_B_Q4_0_1<=wdata[18-1:0];
stb_B_Q4_0_2<=(lb.waddr==383)&lb.wren;if (stb_B_Q4_0_2) reg_B_Q4_0_2<=wdata[18-1:0];
stb_B_Q4_0_3<=(lb.waddr==384)&lb.wren;if (stb_B_Q4_0_3) reg_B_Q4_0_3<=wdata[18-1:0];
stb_B_Q4_0_4<=(lb.waddr==385)&lb.wren;if (stb_B_Q4_0_4) reg_B_Q4_0_4<=wdata[18-1:0];
stb_B_Q4_0_5<=(lb.waddr==386)&lb.wren;if (stb_B_Q4_0_5) reg_B_Q4_0_5<=wdata[18-1:0];
stb_B_Q4_0_6<=(lb.waddr==387)&lb.wren;if (stb_B_Q4_0_6) reg_B_Q4_0_6<=wdata[18-1:0];
stb_B_Q4_0_7<=(lb.waddr==388)&lb.wren;if (stb_B_Q4_0_7) reg_B_Q4_0_7<=wdata[18-1:0];
stb_B_Q4_1_0<=(lb.waddr==389)&lb.wren;if (stb_B_Q4_1_0) reg_B_Q4_1_0<=wdata[18-1:0];
stb_B_Q4_1_1<=(lb.waddr==390)&lb.wren;if (stb_B_Q4_1_1) reg_B_Q4_1_1<=wdata[18-1:0];
stb_B_Q4_1_2<=(lb.waddr==391)&lb.wren;if (stb_B_Q4_1_2) reg_B_Q4_1_2<=wdata[18-1:0];
stb_B_Q4_1_3<=(lb.waddr==392)&lb.wren;if (stb_B_Q4_1_3) reg_B_Q4_1_3<=wdata[18-1:0];
stb_B_Q4_2_0<=(lb.waddr==393)&lb.wren;if (stb_B_Q4_2_0) reg_B_Q4_2_0<=wdata[18-1:0];
stb_W_Q5_0_0_0<=(lb.waddr==394)&lb.wren;if (stb_W_Q5_0_0_0) reg_W_Q5_0_0_0<=wdata[18-1:0];
stb_W_Q5_0_0_1<=(lb.waddr==395)&lb.wren;if (stb_W_Q5_0_0_1) reg_W_Q5_0_0_1<=wdata[18-1:0];
stb_W_Q5_0_0_2<=(lb.waddr==396)&lb.wren;if (stb_W_Q5_0_0_2) reg_W_Q5_0_0_2<=wdata[18-1:0];
stb_W_Q5_0_0_3<=(lb.waddr==397)&lb.wren;if (stb_W_Q5_0_0_3) reg_W_Q5_0_0_3<=wdata[18-1:0];
stb_W_Q5_0_0_4<=(lb.waddr==398)&lb.wren;if (stb_W_Q5_0_0_4) reg_W_Q5_0_0_4<=wdata[18-1:0];
stb_W_Q5_0_0_5<=(lb.waddr==399)&lb.wren;if (stb_W_Q5_0_0_5) reg_W_Q5_0_0_5<=wdata[18-1:0];
stb_W_Q5_0_0_6<=(lb.waddr==400)&lb.wren;if (stb_W_Q5_0_0_6) reg_W_Q5_0_0_6<=wdata[18-1:0];
stb_W_Q5_0_0_7<=(lb.waddr==401)&lb.wren;if (stb_W_Q5_0_0_7) reg_W_Q5_0_0_7<=wdata[18-1:0];
stb_W_Q5_0_1_0<=(lb.waddr==402)&lb.wren;if (stb_W_Q5_0_1_0) reg_W_Q5_0_1_0<=wdata[18-1:0];
stb_W_Q5_0_1_1<=(lb.waddr==403)&lb.wren;if (stb_W_Q5_0_1_1) reg_W_Q5_0_1_1<=wdata[18-1:0];
stb_W_Q5_0_1_2<=(lb.waddr==404)&lb.wren;if (stb_W_Q5_0_1_2) reg_W_Q5_0_1_2<=wdata[18-1:0];
stb_W_Q5_0_1_3<=(lb.waddr==405)&lb.wren;if (stb_W_Q5_0_1_3) reg_W_Q5_0_1_3<=wdata[18-1:0];
stb_W_Q5_0_1_4<=(lb.waddr==406)&lb.wren;if (stb_W_Q5_0_1_4) reg_W_Q5_0_1_4<=wdata[18-1:0];
stb_W_Q5_0_1_5<=(lb.waddr==407)&lb.wren;if (stb_W_Q5_0_1_5) reg_W_Q5_0_1_5<=wdata[18-1:0];
stb_W_Q5_0_1_6<=(lb.waddr==408)&lb.wren;if (stb_W_Q5_0_1_6) reg_W_Q5_0_1_6<=wdata[18-1:0];
stb_W_Q5_0_1_7<=(lb.waddr==409)&lb.wren;if (stb_W_Q5_0_1_7) reg_W_Q5_0_1_7<=wdata[18-1:0];
stb_W_Q5_1_0_0<=(lb.waddr==410)&lb.wren;if (stb_W_Q5_1_0_0) reg_W_Q5_1_0_0<=wdata[18-1:0];
stb_W_Q5_1_0_1<=(lb.waddr==411)&lb.wren;if (stb_W_Q5_1_0_1) reg_W_Q5_1_0_1<=wdata[18-1:0];
stb_W_Q5_1_0_2<=(lb.waddr==412)&lb.wren;if (stb_W_Q5_1_0_2) reg_W_Q5_1_0_2<=wdata[18-1:0];
stb_W_Q5_1_0_3<=(lb.waddr==413)&lb.wren;if (stb_W_Q5_1_0_3) reg_W_Q5_1_0_3<=wdata[18-1:0];
stb_W_Q5_1_1_0<=(lb.waddr==414)&lb.wren;if (stb_W_Q5_1_1_0) reg_W_Q5_1_1_0<=wdata[18-1:0];
stb_W_Q5_1_1_1<=(lb.waddr==415)&lb.wren;if (stb_W_Q5_1_1_1) reg_W_Q5_1_1_1<=wdata[18-1:0];
stb_W_Q5_1_1_2<=(lb.waddr==416)&lb.wren;if (stb_W_Q5_1_1_2) reg_W_Q5_1_1_2<=wdata[18-1:0];
stb_W_Q5_1_1_3<=(lb.waddr==417)&lb.wren;if (stb_W_Q5_1_1_3) reg_W_Q5_1_1_3<=wdata[18-1:0];
stb_W_Q5_1_2_0<=(lb.waddr==418)&lb.wren;if (stb_W_Q5_1_2_0) reg_W_Q5_1_2_0<=wdata[18-1:0];
stb_W_Q5_1_2_1<=(lb.waddr==419)&lb.wren;if (stb_W_Q5_1_2_1) reg_W_Q5_1_2_1<=wdata[18-1:0];
stb_W_Q5_1_2_2<=(lb.waddr==420)&lb.wren;if (stb_W_Q5_1_2_2) reg_W_Q5_1_2_2<=wdata[18-1:0];
stb_W_Q5_1_2_3<=(lb.waddr==421)&lb.wren;if (stb_W_Q5_1_2_3) reg_W_Q5_1_2_3<=wdata[18-1:0];
stb_W_Q5_1_3_0<=(lb.waddr==422)&lb.wren;if (stb_W_Q5_1_3_0) reg_W_Q5_1_3_0<=wdata[18-1:0];
stb_W_Q5_1_3_1<=(lb.waddr==423)&lb.wren;if (stb_W_Q5_1_3_1) reg_W_Q5_1_3_1<=wdata[18-1:0];
stb_W_Q5_1_3_2<=(lb.waddr==424)&lb.wren;if (stb_W_Q5_1_3_2) reg_W_Q5_1_3_2<=wdata[18-1:0];
stb_W_Q5_1_3_3<=(lb.waddr==425)&lb.wren;if (stb_W_Q5_1_3_3) reg_W_Q5_1_3_3<=wdata[18-1:0];
stb_W_Q5_1_4_0<=(lb.waddr==426)&lb.wren;if (stb_W_Q5_1_4_0) reg_W_Q5_1_4_0<=wdata[18-1:0];
stb_W_Q5_1_4_1<=(lb.waddr==427)&lb.wren;if (stb_W_Q5_1_4_1) reg_W_Q5_1_4_1<=wdata[18-1:0];
stb_W_Q5_1_4_2<=(lb.waddr==428)&lb.wren;if (stb_W_Q5_1_4_2) reg_W_Q5_1_4_2<=wdata[18-1:0];
stb_W_Q5_1_4_3<=(lb.waddr==429)&lb.wren;if (stb_W_Q5_1_4_3) reg_W_Q5_1_4_3<=wdata[18-1:0];
stb_W_Q5_1_5_0<=(lb.waddr==430)&lb.wren;if (stb_W_Q5_1_5_0) reg_W_Q5_1_5_0<=wdata[18-1:0];
stb_W_Q5_1_5_1<=(lb.waddr==431)&lb.wren;if (stb_W_Q5_1_5_1) reg_W_Q5_1_5_1<=wdata[18-1:0];
stb_W_Q5_1_5_2<=(lb.waddr==432)&lb.wren;if (stb_W_Q5_1_5_2) reg_W_Q5_1_5_2<=wdata[18-1:0];
stb_W_Q5_1_5_3<=(lb.waddr==433)&lb.wren;if (stb_W_Q5_1_5_3) reg_W_Q5_1_5_3<=wdata[18-1:0];
stb_W_Q5_1_6_0<=(lb.waddr==434)&lb.wren;if (stb_W_Q5_1_6_0) reg_W_Q5_1_6_0<=wdata[18-1:0];
stb_W_Q5_1_6_1<=(lb.waddr==435)&lb.wren;if (stb_W_Q5_1_6_1) reg_W_Q5_1_6_1<=wdata[18-1:0];
stb_W_Q5_1_6_2<=(lb.waddr==436)&lb.wren;if (stb_W_Q5_1_6_2) reg_W_Q5_1_6_2<=wdata[18-1:0];
stb_W_Q5_1_6_3<=(lb.waddr==437)&lb.wren;if (stb_W_Q5_1_6_3) reg_W_Q5_1_6_3<=wdata[18-1:0];
stb_W_Q5_1_7_0<=(lb.waddr==438)&lb.wren;if (stb_W_Q5_1_7_0) reg_W_Q5_1_7_0<=wdata[18-1:0];
stb_W_Q5_1_7_1<=(lb.waddr==439)&lb.wren;if (stb_W_Q5_1_7_1) reg_W_Q5_1_7_1<=wdata[18-1:0];
stb_W_Q5_1_7_2<=(lb.waddr==440)&lb.wren;if (stb_W_Q5_1_7_2) reg_W_Q5_1_7_2<=wdata[18-1:0];
stb_W_Q5_1_7_3<=(lb.waddr==441)&lb.wren;if (stb_W_Q5_1_7_3) reg_W_Q5_1_7_3<=wdata[18-1:0];
stb_W_Q5_2_0_0<=(lb.waddr==442)&lb.wren;if (stb_W_Q5_2_0_0) reg_W_Q5_2_0_0<=wdata[18-1:0];
stb_W_Q5_2_1_0<=(lb.waddr==443)&lb.wren;if (stb_W_Q5_2_1_0) reg_W_Q5_2_1_0<=wdata[18-1:0];
stb_W_Q5_2_2_0<=(lb.waddr==444)&lb.wren;if (stb_W_Q5_2_2_0) reg_W_Q5_2_2_0<=wdata[18-1:0];
stb_W_Q5_2_3_0<=(lb.waddr==445)&lb.wren;if (stb_W_Q5_2_3_0) reg_W_Q5_2_3_0<=wdata[18-1:0];
stb_B_Q5_0_0<=(lb.waddr==446)&lb.wren;if (stb_B_Q5_0_0) reg_B_Q5_0_0<=wdata[18-1:0];
stb_B_Q5_0_1<=(lb.waddr==447)&lb.wren;if (stb_B_Q5_0_1) reg_B_Q5_0_1<=wdata[18-1:0];
stb_B_Q5_0_2<=(lb.waddr==448)&lb.wren;if (stb_B_Q5_0_2) reg_B_Q5_0_2<=wdata[18-1:0];
stb_B_Q5_0_3<=(lb.waddr==449)&lb.wren;if (stb_B_Q5_0_3) reg_B_Q5_0_3<=wdata[18-1:0];
stb_B_Q5_0_4<=(lb.waddr==450)&lb.wren;if (stb_B_Q5_0_4) reg_B_Q5_0_4<=wdata[18-1:0];
stb_B_Q5_0_5<=(lb.waddr==451)&lb.wren;if (stb_B_Q5_0_5) reg_B_Q5_0_5<=wdata[18-1:0];
stb_B_Q5_0_6<=(lb.waddr==452)&lb.wren;if (stb_B_Q5_0_6) reg_B_Q5_0_6<=wdata[18-1:0];
stb_B_Q5_0_7<=(lb.waddr==453)&lb.wren;if (stb_B_Q5_0_7) reg_B_Q5_0_7<=wdata[18-1:0];
stb_B_Q5_1_0<=(lb.waddr==454)&lb.wren;if (stb_B_Q5_1_0) reg_B_Q5_1_0<=wdata[18-1:0];
stb_B_Q5_1_1<=(lb.waddr==455)&lb.wren;if (stb_B_Q5_1_1) reg_B_Q5_1_1<=wdata[18-1:0];
stb_B_Q5_1_2<=(lb.waddr==456)&lb.wren;if (stb_B_Q5_1_2) reg_B_Q5_1_2<=wdata[18-1:0];
stb_B_Q5_1_3<=(lb.waddr==457)&lb.wren;if (stb_B_Q5_1_3) reg_B_Q5_1_3<=wdata[18-1:0];
stb_B_Q5_2_0<=(lb.waddr==458)&lb.wren;if (stb_B_Q5_2_0) reg_B_Q5_2_0<=wdata[18-1:0];
stb_W_Q6_0_0_0<=(lb.waddr==459)&lb.wren;if (stb_W_Q6_0_0_0) reg_W_Q6_0_0_0<=wdata[18-1:0];
stb_W_Q6_0_0_1<=(lb.waddr==460)&lb.wren;if (stb_W_Q6_0_0_1) reg_W_Q6_0_0_1<=wdata[18-1:0];
stb_W_Q6_0_0_2<=(lb.waddr==461)&lb.wren;if (stb_W_Q6_0_0_2) reg_W_Q6_0_0_2<=wdata[18-1:0];
stb_W_Q6_0_0_3<=(lb.waddr==462)&lb.wren;if (stb_W_Q6_0_0_3) reg_W_Q6_0_0_3<=wdata[18-1:0];
stb_W_Q6_0_0_4<=(lb.waddr==463)&lb.wren;if (stb_W_Q6_0_0_4) reg_W_Q6_0_0_4<=wdata[18-1:0];
stb_W_Q6_0_0_5<=(lb.waddr==464)&lb.wren;if (stb_W_Q6_0_0_5) reg_W_Q6_0_0_5<=wdata[18-1:0];
stb_W_Q6_0_0_6<=(lb.waddr==465)&lb.wren;if (stb_W_Q6_0_0_6) reg_W_Q6_0_0_6<=wdata[18-1:0];
stb_W_Q6_0_0_7<=(lb.waddr==466)&lb.wren;if (stb_W_Q6_0_0_7) reg_W_Q6_0_0_7<=wdata[18-1:0];
stb_W_Q6_0_1_0<=(lb.waddr==467)&lb.wren;if (stb_W_Q6_0_1_0) reg_W_Q6_0_1_0<=wdata[18-1:0];
stb_W_Q6_0_1_1<=(lb.waddr==468)&lb.wren;if (stb_W_Q6_0_1_1) reg_W_Q6_0_1_1<=wdata[18-1:0];
stb_W_Q6_0_1_2<=(lb.waddr==469)&lb.wren;if (stb_W_Q6_0_1_2) reg_W_Q6_0_1_2<=wdata[18-1:0];
stb_W_Q6_0_1_3<=(lb.waddr==470)&lb.wren;if (stb_W_Q6_0_1_3) reg_W_Q6_0_1_3<=wdata[18-1:0];
stb_W_Q6_0_1_4<=(lb.waddr==471)&lb.wren;if (stb_W_Q6_0_1_4) reg_W_Q6_0_1_4<=wdata[18-1:0];
stb_W_Q6_0_1_5<=(lb.waddr==472)&lb.wren;if (stb_W_Q6_0_1_5) reg_W_Q6_0_1_5<=wdata[18-1:0];
stb_W_Q6_0_1_6<=(lb.waddr==473)&lb.wren;if (stb_W_Q6_0_1_6) reg_W_Q6_0_1_6<=wdata[18-1:0];
stb_W_Q6_0_1_7<=(lb.waddr==474)&lb.wren;if (stb_W_Q6_0_1_7) reg_W_Q6_0_1_7<=wdata[18-1:0];
stb_W_Q6_1_0_0<=(lb.waddr==475)&lb.wren;if (stb_W_Q6_1_0_0) reg_W_Q6_1_0_0<=wdata[18-1:0];
stb_W_Q6_1_0_1<=(lb.waddr==476)&lb.wren;if (stb_W_Q6_1_0_1) reg_W_Q6_1_0_1<=wdata[18-1:0];
stb_W_Q6_1_0_2<=(lb.waddr==477)&lb.wren;if (stb_W_Q6_1_0_2) reg_W_Q6_1_0_2<=wdata[18-1:0];
stb_W_Q6_1_0_3<=(lb.waddr==478)&lb.wren;if (stb_W_Q6_1_0_3) reg_W_Q6_1_0_3<=wdata[18-1:0];
stb_W_Q6_1_1_0<=(lb.waddr==479)&lb.wren;if (stb_W_Q6_1_1_0) reg_W_Q6_1_1_0<=wdata[18-1:0];
stb_W_Q6_1_1_1<=(lb.waddr==480)&lb.wren;if (stb_W_Q6_1_1_1) reg_W_Q6_1_1_1<=wdata[18-1:0];
stb_W_Q6_1_1_2<=(lb.waddr==481)&lb.wren;if (stb_W_Q6_1_1_2) reg_W_Q6_1_1_2<=wdata[18-1:0];
stb_W_Q6_1_1_3<=(lb.waddr==482)&lb.wren;if (stb_W_Q6_1_1_3) reg_W_Q6_1_1_3<=wdata[18-1:0];
stb_W_Q6_1_2_0<=(lb.waddr==483)&lb.wren;if (stb_W_Q6_1_2_0) reg_W_Q6_1_2_0<=wdata[18-1:0];
stb_W_Q6_1_2_1<=(lb.waddr==484)&lb.wren;if (stb_W_Q6_1_2_1) reg_W_Q6_1_2_1<=wdata[18-1:0];
stb_W_Q6_1_2_2<=(lb.waddr==485)&lb.wren;if (stb_W_Q6_1_2_2) reg_W_Q6_1_2_2<=wdata[18-1:0];
stb_W_Q6_1_2_3<=(lb.waddr==486)&lb.wren;if (stb_W_Q6_1_2_3) reg_W_Q6_1_2_3<=wdata[18-1:0];
stb_W_Q6_1_3_0<=(lb.waddr==487)&lb.wren;if (stb_W_Q6_1_3_0) reg_W_Q6_1_3_0<=wdata[18-1:0];
stb_W_Q6_1_3_1<=(lb.waddr==488)&lb.wren;if (stb_W_Q6_1_3_1) reg_W_Q6_1_3_1<=wdata[18-1:0];
stb_W_Q6_1_3_2<=(lb.waddr==489)&lb.wren;if (stb_W_Q6_1_3_2) reg_W_Q6_1_3_2<=wdata[18-1:0];
stb_W_Q6_1_3_3<=(lb.waddr==490)&lb.wren;if (stb_W_Q6_1_3_3) reg_W_Q6_1_3_3<=wdata[18-1:0];
stb_W_Q6_1_4_0<=(lb.waddr==491)&lb.wren;if (stb_W_Q6_1_4_0) reg_W_Q6_1_4_0<=wdata[18-1:0];
stb_W_Q6_1_4_1<=(lb.waddr==492)&lb.wren;if (stb_W_Q6_1_4_1) reg_W_Q6_1_4_1<=wdata[18-1:0];
stb_W_Q6_1_4_2<=(lb.waddr==493)&lb.wren;if (stb_W_Q6_1_4_2) reg_W_Q6_1_4_2<=wdata[18-1:0];
stb_W_Q6_1_4_3<=(lb.waddr==494)&lb.wren;if (stb_W_Q6_1_4_3) reg_W_Q6_1_4_3<=wdata[18-1:0];
stb_W_Q6_1_5_0<=(lb.waddr==495)&lb.wren;if (stb_W_Q6_1_5_0) reg_W_Q6_1_5_0<=wdata[18-1:0];
stb_W_Q6_1_5_1<=(lb.waddr==496)&lb.wren;if (stb_W_Q6_1_5_1) reg_W_Q6_1_5_1<=wdata[18-1:0];
stb_W_Q6_1_5_2<=(lb.waddr==497)&lb.wren;if (stb_W_Q6_1_5_2) reg_W_Q6_1_5_2<=wdata[18-1:0];
stb_W_Q6_1_5_3<=(lb.waddr==498)&lb.wren;if (stb_W_Q6_1_5_3) reg_W_Q6_1_5_3<=wdata[18-1:0];
stb_W_Q6_1_6_0<=(lb.waddr==499)&lb.wren;if (stb_W_Q6_1_6_0) reg_W_Q6_1_6_0<=wdata[18-1:0];
stb_W_Q6_1_6_1<=(lb.waddr==500)&lb.wren;if (stb_W_Q6_1_6_1) reg_W_Q6_1_6_1<=wdata[18-1:0];
stb_W_Q6_1_6_2<=(lb.waddr==501)&lb.wren;if (stb_W_Q6_1_6_2) reg_W_Q6_1_6_2<=wdata[18-1:0];
stb_W_Q6_1_6_3<=(lb.waddr==502)&lb.wren;if (stb_W_Q6_1_6_3) reg_W_Q6_1_6_3<=wdata[18-1:0];
stb_W_Q6_1_7_0<=(lb.waddr==503)&lb.wren;if (stb_W_Q6_1_7_0) reg_W_Q6_1_7_0<=wdata[18-1:0];
stb_W_Q6_1_7_1<=(lb.waddr==504)&lb.wren;if (stb_W_Q6_1_7_1) reg_W_Q6_1_7_1<=wdata[18-1:0];
stb_W_Q6_1_7_2<=(lb.waddr==505)&lb.wren;if (stb_W_Q6_1_7_2) reg_W_Q6_1_7_2<=wdata[18-1:0];
stb_W_Q6_1_7_3<=(lb.waddr==506)&lb.wren;if (stb_W_Q6_1_7_3) reg_W_Q6_1_7_3<=wdata[18-1:0];
stb_W_Q6_2_0_0<=(lb.waddr==507)&lb.wren;if (stb_W_Q6_2_0_0) reg_W_Q6_2_0_0<=wdata[18-1:0];
stb_W_Q6_2_1_0<=(lb.waddr==508)&lb.wren;if (stb_W_Q6_2_1_0) reg_W_Q6_2_1_0<=wdata[18-1:0];
stb_W_Q6_2_2_0<=(lb.waddr==509)&lb.wren;if (stb_W_Q6_2_2_0) reg_W_Q6_2_2_0<=wdata[18-1:0];
stb_W_Q6_2_3_0<=(lb.waddr==510)&lb.wren;if (stb_W_Q6_2_3_0) reg_W_Q6_2_3_0<=wdata[18-1:0];
stb_B_Q6_0_0<=(lb.waddr==511)&lb.wren;if (stb_B_Q6_0_0) reg_B_Q6_0_0<=wdata[18-1:0];
stb_B_Q6_0_1<=(lb.waddr==512)&lb.wren;if (stb_B_Q6_0_1) reg_B_Q6_0_1<=wdata[18-1:0];
stb_B_Q6_0_2<=(lb.waddr==513)&lb.wren;if (stb_B_Q6_0_2) reg_B_Q6_0_2<=wdata[18-1:0];
stb_B_Q6_0_3<=(lb.waddr==514)&lb.wren;if (stb_B_Q6_0_3) reg_B_Q6_0_3<=wdata[18-1:0];
stb_B_Q6_0_4<=(lb.waddr==515)&lb.wren;if (stb_B_Q6_0_4) reg_B_Q6_0_4<=wdata[18-1:0];
stb_B_Q6_0_5<=(lb.waddr==516)&lb.wren;if (stb_B_Q6_0_5) reg_B_Q6_0_5<=wdata[18-1:0];
stb_B_Q6_0_6<=(lb.waddr==517)&lb.wren;if (stb_B_Q6_0_6) reg_B_Q6_0_6<=wdata[18-1:0];
stb_B_Q6_0_7<=(lb.waddr==518)&lb.wren;if (stb_B_Q6_0_7) reg_B_Q6_0_7<=wdata[18-1:0];
stb_B_Q6_1_0<=(lb.waddr==519)&lb.wren;if (stb_B_Q6_1_0) reg_B_Q6_1_0<=wdata[18-1:0];
stb_B_Q6_1_1<=(lb.waddr==520)&lb.wren;if (stb_B_Q6_1_1) reg_B_Q6_1_1<=wdata[18-1:0];
stb_B_Q6_1_2<=(lb.waddr==521)&lb.wren;if (stb_B_Q6_1_2) reg_B_Q6_1_2<=wdata[18-1:0];
stb_B_Q6_1_3<=(lb.waddr==522)&lb.wren;if (stb_B_Q6_1_3) reg_B_Q6_1_3<=wdata[18-1:0];
stb_B_Q6_2_0<=(lb.waddr==523)&lb.wren;if (stb_B_Q6_2_0) reg_B_Q6_2_0<=wdata[18-1:0];
stb_W_Q7_0_0_0<=(lb.waddr==524)&lb.wren;if (stb_W_Q7_0_0_0) reg_W_Q7_0_0_0<=wdata[18-1:0];
stb_W_Q7_0_0_1<=(lb.waddr==525)&lb.wren;if (stb_W_Q7_0_0_1) reg_W_Q7_0_0_1<=wdata[18-1:0];
stb_W_Q7_0_0_2<=(lb.waddr==526)&lb.wren;if (stb_W_Q7_0_0_2) reg_W_Q7_0_0_2<=wdata[18-1:0];
stb_W_Q7_0_0_3<=(lb.waddr==527)&lb.wren;if (stb_W_Q7_0_0_3) reg_W_Q7_0_0_3<=wdata[18-1:0];
stb_W_Q7_0_0_4<=(lb.waddr==528)&lb.wren;if (stb_W_Q7_0_0_4) reg_W_Q7_0_0_4<=wdata[18-1:0];
stb_W_Q7_0_0_5<=(lb.waddr==529)&lb.wren;if (stb_W_Q7_0_0_5) reg_W_Q7_0_0_5<=wdata[18-1:0];
stb_W_Q7_0_0_6<=(lb.waddr==530)&lb.wren;if (stb_W_Q7_0_0_6) reg_W_Q7_0_0_6<=wdata[18-1:0];
stb_W_Q7_0_0_7<=(lb.waddr==531)&lb.wren;if (stb_W_Q7_0_0_7) reg_W_Q7_0_0_7<=wdata[18-1:0];
stb_W_Q7_0_1_0<=(lb.waddr==532)&lb.wren;if (stb_W_Q7_0_1_0) reg_W_Q7_0_1_0<=wdata[18-1:0];
stb_W_Q7_0_1_1<=(lb.waddr==533)&lb.wren;if (stb_W_Q7_0_1_1) reg_W_Q7_0_1_1<=wdata[18-1:0];
stb_W_Q7_0_1_2<=(lb.waddr==534)&lb.wren;if (stb_W_Q7_0_1_2) reg_W_Q7_0_1_2<=wdata[18-1:0];
stb_W_Q7_0_1_3<=(lb.waddr==535)&lb.wren;if (stb_W_Q7_0_1_3) reg_W_Q7_0_1_3<=wdata[18-1:0];
stb_W_Q7_0_1_4<=(lb.waddr==536)&lb.wren;if (stb_W_Q7_0_1_4) reg_W_Q7_0_1_4<=wdata[18-1:0];
stb_W_Q7_0_1_5<=(lb.waddr==537)&lb.wren;if (stb_W_Q7_0_1_5) reg_W_Q7_0_1_5<=wdata[18-1:0];
stb_W_Q7_0_1_6<=(lb.waddr==538)&lb.wren;if (stb_W_Q7_0_1_6) reg_W_Q7_0_1_6<=wdata[18-1:0];
stb_W_Q7_0_1_7<=(lb.waddr==539)&lb.wren;if (stb_W_Q7_0_1_7) reg_W_Q7_0_1_7<=wdata[18-1:0];
stb_W_Q7_1_0_0<=(lb.waddr==540)&lb.wren;if (stb_W_Q7_1_0_0) reg_W_Q7_1_0_0<=wdata[18-1:0];
stb_W_Q7_1_0_1<=(lb.waddr==541)&lb.wren;if (stb_W_Q7_1_0_1) reg_W_Q7_1_0_1<=wdata[18-1:0];
stb_W_Q7_1_0_2<=(lb.waddr==542)&lb.wren;if (stb_W_Q7_1_0_2) reg_W_Q7_1_0_2<=wdata[18-1:0];
stb_W_Q7_1_0_3<=(lb.waddr==543)&lb.wren;if (stb_W_Q7_1_0_3) reg_W_Q7_1_0_3<=wdata[18-1:0];
stb_W_Q7_1_1_0<=(lb.waddr==544)&lb.wren;if (stb_W_Q7_1_1_0) reg_W_Q7_1_1_0<=wdata[18-1:0];
stb_W_Q7_1_1_1<=(lb.waddr==545)&lb.wren;if (stb_W_Q7_1_1_1) reg_W_Q7_1_1_1<=wdata[18-1:0];
stb_W_Q7_1_1_2<=(lb.waddr==546)&lb.wren;if (stb_W_Q7_1_1_2) reg_W_Q7_1_1_2<=wdata[18-1:0];
stb_W_Q7_1_1_3<=(lb.waddr==547)&lb.wren;if (stb_W_Q7_1_1_3) reg_W_Q7_1_1_3<=wdata[18-1:0];
stb_W_Q7_1_2_0<=(lb.waddr==548)&lb.wren;if (stb_W_Q7_1_2_0) reg_W_Q7_1_2_0<=wdata[18-1:0];
stb_W_Q7_1_2_1<=(lb.waddr==549)&lb.wren;if (stb_W_Q7_1_2_1) reg_W_Q7_1_2_1<=wdata[18-1:0];
stb_W_Q7_1_2_2<=(lb.waddr==550)&lb.wren;if (stb_W_Q7_1_2_2) reg_W_Q7_1_2_2<=wdata[18-1:0];
stb_W_Q7_1_2_3<=(lb.waddr==551)&lb.wren;if (stb_W_Q7_1_2_3) reg_W_Q7_1_2_3<=wdata[18-1:0];
stb_W_Q7_1_3_0<=(lb.waddr==552)&lb.wren;if (stb_W_Q7_1_3_0) reg_W_Q7_1_3_0<=wdata[18-1:0];
stb_W_Q7_1_3_1<=(lb.waddr==553)&lb.wren;if (stb_W_Q7_1_3_1) reg_W_Q7_1_3_1<=wdata[18-1:0];
stb_W_Q7_1_3_2<=(lb.waddr==554)&lb.wren;if (stb_W_Q7_1_3_2) reg_W_Q7_1_3_2<=wdata[18-1:0];
stb_W_Q7_1_3_3<=(lb.waddr==555)&lb.wren;if (stb_W_Q7_1_3_3) reg_W_Q7_1_3_3<=wdata[18-1:0];
stb_W_Q7_1_4_0<=(lb.waddr==556)&lb.wren;if (stb_W_Q7_1_4_0) reg_W_Q7_1_4_0<=wdata[18-1:0];
stb_W_Q7_1_4_1<=(lb.waddr==557)&lb.wren;if (stb_W_Q7_1_4_1) reg_W_Q7_1_4_1<=wdata[18-1:0];
stb_W_Q7_1_4_2<=(lb.waddr==558)&lb.wren;if (stb_W_Q7_1_4_2) reg_W_Q7_1_4_2<=wdata[18-1:0];
stb_W_Q7_1_4_3<=(lb.waddr==559)&lb.wren;if (stb_W_Q7_1_4_3) reg_W_Q7_1_4_3<=wdata[18-1:0];
stb_W_Q7_1_5_0<=(lb.waddr==560)&lb.wren;if (stb_W_Q7_1_5_0) reg_W_Q7_1_5_0<=wdata[18-1:0];
stb_W_Q7_1_5_1<=(lb.waddr==561)&lb.wren;if (stb_W_Q7_1_5_1) reg_W_Q7_1_5_1<=wdata[18-1:0];
stb_W_Q7_1_5_2<=(lb.waddr==562)&lb.wren;if (stb_W_Q7_1_5_2) reg_W_Q7_1_5_2<=wdata[18-1:0];
stb_W_Q7_1_5_3<=(lb.waddr==563)&lb.wren;if (stb_W_Q7_1_5_3) reg_W_Q7_1_5_3<=wdata[18-1:0];
stb_W_Q7_1_6_0<=(lb.waddr==564)&lb.wren;if (stb_W_Q7_1_6_0) reg_W_Q7_1_6_0<=wdata[18-1:0];
stb_W_Q7_1_6_1<=(lb.waddr==565)&lb.wren;if (stb_W_Q7_1_6_1) reg_W_Q7_1_6_1<=wdata[18-1:0];
stb_W_Q7_1_6_2<=(lb.waddr==566)&lb.wren;if (stb_W_Q7_1_6_2) reg_W_Q7_1_6_2<=wdata[18-1:0];
stb_W_Q7_1_6_3<=(lb.waddr==567)&lb.wren;if (stb_W_Q7_1_6_3) reg_W_Q7_1_6_3<=wdata[18-1:0];
stb_W_Q7_1_7_0<=(lb.waddr==568)&lb.wren;if (stb_W_Q7_1_7_0) reg_W_Q7_1_7_0<=wdata[18-1:0];
stb_W_Q7_1_7_1<=(lb.waddr==569)&lb.wren;if (stb_W_Q7_1_7_1) reg_W_Q7_1_7_1<=wdata[18-1:0];
stb_W_Q7_1_7_2<=(lb.waddr==570)&lb.wren;if (stb_W_Q7_1_7_2) reg_W_Q7_1_7_2<=wdata[18-1:0];
stb_W_Q7_1_7_3<=(lb.waddr==571)&lb.wren;if (stb_W_Q7_1_7_3) reg_W_Q7_1_7_3<=wdata[18-1:0];
stb_W_Q7_2_0_0<=(lb.waddr==572)&lb.wren;if (stb_W_Q7_2_0_0) reg_W_Q7_2_0_0<=wdata[18-1:0];
stb_W_Q7_2_1_0<=(lb.waddr==573)&lb.wren;if (stb_W_Q7_2_1_0) reg_W_Q7_2_1_0<=wdata[18-1:0];
stb_W_Q7_2_2_0<=(lb.waddr==574)&lb.wren;if (stb_W_Q7_2_2_0) reg_W_Q7_2_2_0<=wdata[18-1:0];
stb_W_Q7_2_3_0<=(lb.waddr==575)&lb.wren;if (stb_W_Q7_2_3_0) reg_W_Q7_2_3_0<=wdata[18-1:0];
stb_B_Q7_0_0<=(lb.waddr==576)&lb.wren;if (stb_B_Q7_0_0) reg_B_Q7_0_0<=wdata[18-1:0];
stb_B_Q7_0_1<=(lb.waddr==577)&lb.wren;if (stb_B_Q7_0_1) reg_B_Q7_0_1<=wdata[18-1:0];
stb_B_Q7_0_2<=(lb.waddr==578)&lb.wren;if (stb_B_Q7_0_2) reg_B_Q7_0_2<=wdata[18-1:0];
stb_B_Q7_0_3<=(lb.waddr==579)&lb.wren;if (stb_B_Q7_0_3) reg_B_Q7_0_3<=wdata[18-1:0];
stb_B_Q7_0_4<=(lb.waddr==580)&lb.wren;if (stb_B_Q7_0_4) reg_B_Q7_0_4<=wdata[18-1:0];
stb_B_Q7_0_5<=(lb.waddr==581)&lb.wren;if (stb_B_Q7_0_5) reg_B_Q7_0_5<=wdata[18-1:0];
stb_B_Q7_0_6<=(lb.waddr==582)&lb.wren;if (stb_B_Q7_0_6) reg_B_Q7_0_6<=wdata[18-1:0];
stb_B_Q7_0_7<=(lb.waddr==583)&lb.wren;if (stb_B_Q7_0_7) reg_B_Q7_0_7<=wdata[18-1:0];
stb_B_Q7_1_0<=(lb.waddr==584)&lb.wren;if (stb_B_Q7_1_0) reg_B_Q7_1_0<=wdata[18-1:0];
stb_B_Q7_1_1<=(lb.waddr==585)&lb.wren;if (stb_B_Q7_1_1) reg_B_Q7_1_1<=wdata[18-1:0];
stb_B_Q7_1_2<=(lb.waddr==586)&lb.wren;if (stb_B_Q7_1_2) reg_B_Q7_1_2<=wdata[18-1:0];
stb_B_Q7_1_3<=(lb.waddr==587)&lb.wren;if (stb_B_Q7_1_3) reg_B_Q7_1_3<=wdata[18-1:0];
stb_B_Q7_2_0<=(lb.waddr==588)&lb.wren;if (stb_B_Q7_2_0) reg_B_Q7_2_0<=wdata[18-1:0];
stb_min_Q0_I<=(lb.waddr==589)&lb.wren;if (stb_min_Q0_I) reg_min_Q0_I<=wdata[32-1:0];
stb_min_Q0_Q<=(lb.waddr==590)&lb.wren;if (stb_min_Q0_Q) reg_min_Q0_Q<=wdata[32-1:0];
stb_min_Q1_I<=(lb.waddr==591)&lb.wren;if (stb_min_Q1_I) reg_min_Q1_I<=wdata[32-1:0];
stb_min_Q1_Q<=(lb.waddr==592)&lb.wren;if (stb_min_Q1_Q) reg_min_Q1_Q<=wdata[32-1:0];
stb_min_Q2_I<=(lb.waddr==593)&lb.wren;if (stb_min_Q2_I) reg_min_Q2_I<=wdata[32-1:0];
stb_min_Q2_Q<=(lb.waddr==594)&lb.wren;if (stb_min_Q2_Q) reg_min_Q2_Q<=wdata[32-1:0];
stb_min_Q3_I<=(lb.waddr==595)&lb.wren;if (stb_min_Q3_I) reg_min_Q3_I<=wdata[32-1:0];
stb_min_Q3_Q<=(lb.waddr==596)&lb.wren;if (stb_min_Q3_Q) reg_min_Q3_Q<=wdata[32-1:0];
stb_min_Q4_I<=(lb.waddr==597)&lb.wren;if (stb_min_Q4_I) reg_min_Q4_I<=wdata[32-1:0];
stb_min_Q4_Q<=(lb.waddr==598)&lb.wren;if (stb_min_Q4_Q) reg_min_Q4_Q<=wdata[32-1:0];
stb_min_Q5_I<=(lb.waddr==599)&lb.wren;if (stb_min_Q5_I) reg_min_Q5_I<=wdata[32-1:0];
stb_min_Q5_Q<=(lb.waddr==600)&lb.wren;if (stb_min_Q5_Q) reg_min_Q5_Q<=wdata[32-1:0];
stb_min_Q6_I<=(lb.waddr==601)&lb.wren;if (stb_min_Q6_I) reg_min_Q6_I<=wdata[32-1:0];
stb_min_Q6_Q<=(lb.waddr==602)&lb.wren;if (stb_min_Q6_Q) reg_min_Q6_Q<=wdata[32-1:0];
stb_min_Q7_I<=(lb.waddr==603)&lb.wren;if (stb_min_Q7_I) reg_min_Q7_I<=wdata[32-1:0];
stb_min_Q7_Q<=(lb.waddr==604)&lb.wren;if (stb_min_Q7_Q) reg_min_Q7_Q<=wdata[32-1:0];
end
always @(posedge lb.clk) begin
if (lb.rden16[READDELAY]) begin
case (lb.raddr16[(READDELAY+1)*ADDR_WIDTH-1:READDELAY*ADDR_WIDTH]) 

1: rdata <= resetacc;
2: rdata <= addr_accbuf_mon0;
3: rdata <= addr_accbuf_mon1;
4: rdata <= addr_accbuf_mon2;
5: rdata <= addr_accbuf_mon3;
6: rdata <= amp;
7: rdata <= bramsel;
8: rdata <= busy;
9: rdata <= coef00;
10: rdata <= coef01;
11: rdata <= coef02;
12: rdata <= coef03;
13: rdata <= coef10;
14: rdata <= coef11;
15: rdata <= coef12;
16: rdata <= coef13;
17: rdata <= coef20;
18: rdata <= coef21;
19: rdata <= coef22;
20: rdata <= coef23;
21: rdata <= coef30;
22: rdata <= coef31;
23: rdata <= coef32;
24: rdata <= coef33;
25: rdata <= dacsel;
26: rdata <= dspreset;
27: rdata <= lastshotdone;
28: rdata <= nshot;
29: rdata <= qdrvfreqsel;
30: rdata <= rdlofreqsel;
31: rdata <= rdrvfreqsel;
32: rdata <= reset_bram_read;
33: rdata <= shotcnt;
34: rdata <= start;
35: rdata <= test;
36: rdata <= test1;
37: rdata <= acqbufreset;
38: rdata <= dacmonreset;
39: rdata <= decimator;
40: rdata <= acqchansel0;
41: rdata <= acqchansel1;
42: rdata <= dacmonchansel0;
43: rdata <= dacmonchansel1;
44: rdata <= dacmonchansel2;
45: rdata <= dacmonchansel3;
46: rdata <= delayaftertrig;
47: rdata <= mixbb1sel;
48: rdata <= mixbb2sel;
49: rdata <= shift;
50: rdata <= procdone;
51: rdata <= cnt00;
52: rdata <= cnt01;
53: rdata <= cnt02;
54: rdata <= cnt03;
55: rdata <= cnt10;
56: rdata <= cnt11;
57: rdata <= cnt12;
58: rdata <= cnt13;
59: rdata <= cnt20;
60: rdata <= cnt21;
61: rdata <= cnt22;
62: rdata <= cnt23;
63: rdata <= cnt30;
64: rdata <= cnt31;
65: rdata <= cnt32;
66: rdata <= cnt33;
67: rdata <= addr_sdbuf_mon0;
68: rdata <= addr_sdbuf_mon1;
69: rdata <= W_Q0_0_0_0;
70: rdata <= W_Q0_0_0_1;
71: rdata <= W_Q0_0_0_2;
72: rdata <= W_Q0_0_0_3;
73: rdata <= W_Q0_0_0_4;
74: rdata <= W_Q0_0_0_5;
75: rdata <= W_Q0_0_0_6;
76: rdata <= W_Q0_0_0_7;
77: rdata <= W_Q0_0_1_0;
78: rdata <= W_Q0_0_1_1;
79: rdata <= W_Q0_0_1_2;
80: rdata <= W_Q0_0_1_3;
81: rdata <= W_Q0_0_1_4;
82: rdata <= W_Q0_0_1_5;
83: rdata <= W_Q0_0_1_6;
84: rdata <= W_Q0_0_1_7;
85: rdata <= W_Q0_1_0_0;
86: rdata <= W_Q0_1_0_1;
87: rdata <= W_Q0_1_0_2;
88: rdata <= W_Q0_1_0_3;
89: rdata <= W_Q0_1_1_0;
90: rdata <= W_Q0_1_1_1;
91: rdata <= W_Q0_1_1_2;
92: rdata <= W_Q0_1_1_3;
93: rdata <= W_Q0_1_2_0;
94: rdata <= W_Q0_1_2_1;
95: rdata <= W_Q0_1_2_2;
96: rdata <= W_Q0_1_2_3;
97: rdata <= W_Q0_1_3_0;
98: rdata <= W_Q0_1_3_1;
99: rdata <= W_Q0_1_3_2;
100: rdata <= W_Q0_1_3_3;
101: rdata <= W_Q0_1_4_0;
102: rdata <= W_Q0_1_4_1;
103: rdata <= W_Q0_1_4_2;
104: rdata <= W_Q0_1_4_3;
105: rdata <= W_Q0_1_5_0;
106: rdata <= W_Q0_1_5_1;
107: rdata <= W_Q0_1_5_2;
108: rdata <= W_Q0_1_5_3;
109: rdata <= W_Q0_1_6_0;
110: rdata <= W_Q0_1_6_1;
111: rdata <= W_Q0_1_6_2;
112: rdata <= W_Q0_1_6_3;
113: rdata <= W_Q0_1_7_0;
114: rdata <= W_Q0_1_7_1;
115: rdata <= W_Q0_1_7_2;
116: rdata <= W_Q0_1_7_3;
117: rdata <= W_Q0_2_0_0;
118: rdata <= W_Q0_2_1_0;
119: rdata <= W_Q0_2_2_0;
120: rdata <= W_Q0_2_3_0;
121: rdata <= B_Q0_0_0;
122: rdata <= B_Q0_0_1;
123: rdata <= B_Q0_0_2;
124: rdata <= B_Q0_0_3;
125: rdata <= B_Q0_0_4;
126: rdata <= B_Q0_0_5;
127: rdata <= B_Q0_0_6;
128: rdata <= B_Q0_0_7;
129: rdata <= B_Q0_1_0;
130: rdata <= B_Q0_1_1;
131: rdata <= B_Q0_1_2;
132: rdata <= B_Q0_1_3;
133: rdata <= B_Q0_2_0;
134: rdata <= W_Q1_0_0_0;
135: rdata <= W_Q1_0_0_1;
136: rdata <= W_Q1_0_0_2;
137: rdata <= W_Q1_0_0_3;
138: rdata <= W_Q1_0_0_4;
139: rdata <= W_Q1_0_0_5;
140: rdata <= W_Q1_0_0_6;
141: rdata <= W_Q1_0_0_7;
142: rdata <= W_Q1_0_1_0;
143: rdata <= W_Q1_0_1_1;
144: rdata <= W_Q1_0_1_2;
145: rdata <= W_Q1_0_1_3;
146: rdata <= W_Q1_0_1_4;
147: rdata <= W_Q1_0_1_5;
148: rdata <= W_Q1_0_1_6;
149: rdata <= W_Q1_0_1_7;
150: rdata <= W_Q1_1_0_0;
151: rdata <= W_Q1_1_0_1;
152: rdata <= W_Q1_1_0_2;
153: rdata <= W_Q1_1_0_3;
154: rdata <= W_Q1_1_1_0;
155: rdata <= W_Q1_1_1_1;
156: rdata <= W_Q1_1_1_2;
157: rdata <= W_Q1_1_1_3;
158: rdata <= W_Q1_1_2_0;
159: rdata <= W_Q1_1_2_1;
160: rdata <= W_Q1_1_2_2;
161: rdata <= W_Q1_1_2_3;
162: rdata <= W_Q1_1_3_0;
163: rdata <= W_Q1_1_3_1;
164: rdata <= W_Q1_1_3_2;
165: rdata <= W_Q1_1_3_3;
166: rdata <= W_Q1_1_4_0;
167: rdata <= W_Q1_1_4_1;
168: rdata <= W_Q1_1_4_2;
169: rdata <= W_Q1_1_4_3;
170: rdata <= W_Q1_1_5_0;
171: rdata <= W_Q1_1_5_1;
172: rdata <= W_Q1_1_5_2;
173: rdata <= W_Q1_1_5_3;
174: rdata <= W_Q1_1_6_0;
175: rdata <= W_Q1_1_6_1;
176: rdata <= W_Q1_1_6_2;
177: rdata <= W_Q1_1_6_3;
178: rdata <= W_Q1_1_7_0;
179: rdata <= W_Q1_1_7_1;
180: rdata <= W_Q1_1_7_2;
181: rdata <= W_Q1_1_7_3;
182: rdata <= W_Q1_2_0_0;
183: rdata <= W_Q1_2_1_0;
184: rdata <= W_Q1_2_2_0;
185: rdata <= W_Q1_2_3_0;
186: rdata <= B_Q1_0_0;
187: rdata <= B_Q1_0_1;
188: rdata <= B_Q1_0_2;
189: rdata <= B_Q1_0_3;
190: rdata <= B_Q1_0_4;
191: rdata <= B_Q1_0_5;
192: rdata <= B_Q1_0_6;
193: rdata <= B_Q1_0_7;
194: rdata <= B_Q1_1_0;
195: rdata <= B_Q1_1_1;
196: rdata <= B_Q1_1_2;
197: rdata <= B_Q1_1_3;
198: rdata <= B_Q1_2_0;
199: rdata <= W_Q2_0_0_0;
200: rdata <= W_Q2_0_0_1;
201: rdata <= W_Q2_0_0_2;
202: rdata <= W_Q2_0_0_3;
203: rdata <= W_Q2_0_0_4;
204: rdata <= W_Q2_0_0_5;
205: rdata <= W_Q2_0_0_6;
206: rdata <= W_Q2_0_0_7;
207: rdata <= W_Q2_0_1_0;
208: rdata <= W_Q2_0_1_1;
209: rdata <= W_Q2_0_1_2;
210: rdata <= W_Q2_0_1_3;
211: rdata <= W_Q2_0_1_4;
212: rdata <= W_Q2_0_1_5;
213: rdata <= W_Q2_0_1_6;
214: rdata <= W_Q2_0_1_7;
215: rdata <= W_Q2_1_0_0;
216: rdata <= W_Q2_1_0_1;
217: rdata <= W_Q2_1_0_2;
218: rdata <= W_Q2_1_0_3;
219: rdata <= W_Q2_1_1_0;
220: rdata <= W_Q2_1_1_1;
221: rdata <= W_Q2_1_1_2;
222: rdata <= W_Q2_1_1_3;
223: rdata <= W_Q2_1_2_0;
224: rdata <= W_Q2_1_2_1;
225: rdata <= W_Q2_1_2_2;
226: rdata <= W_Q2_1_2_3;
227: rdata <= W_Q2_1_3_0;
228: rdata <= W_Q2_1_3_1;
229: rdata <= W_Q2_1_3_2;
230: rdata <= W_Q2_1_3_3;
231: rdata <= W_Q2_1_4_0;
232: rdata <= W_Q2_1_4_1;
233: rdata <= W_Q2_1_4_2;
234: rdata <= W_Q2_1_4_3;
235: rdata <= W_Q2_1_5_0;
236: rdata <= W_Q2_1_5_1;
237: rdata <= W_Q2_1_5_2;
238: rdata <= W_Q2_1_5_3;
239: rdata <= W_Q2_1_6_0;
240: rdata <= W_Q2_1_6_1;
241: rdata <= W_Q2_1_6_2;
242: rdata <= W_Q2_1_6_3;
243: rdata <= W_Q2_1_7_0;
244: rdata <= W_Q2_1_7_1;
245: rdata <= W_Q2_1_7_2;
246: rdata <= W_Q2_1_7_3;
247: rdata <= W_Q2_2_0_0;
248: rdata <= W_Q2_2_1_0;
249: rdata <= W_Q2_2_2_0;
250: rdata <= W_Q2_2_3_0;
251: rdata <= B_Q2_0_0;
252: rdata <= B_Q2_0_1;
253: rdata <= B_Q2_0_2;
254: rdata <= B_Q2_0_3;
255: rdata <= B_Q2_0_4;
256: rdata <= B_Q2_0_5;
257: rdata <= B_Q2_0_6;
258: rdata <= B_Q2_0_7;
259: rdata <= B_Q2_1_0;
260: rdata <= B_Q2_1_1;
261: rdata <= B_Q2_1_2;
262: rdata <= B_Q2_1_3;
263: rdata <= B_Q2_2_0;
264: rdata <= W_Q3_0_0_0;
265: rdata <= W_Q3_0_0_1;
266: rdata <= W_Q3_0_0_2;
267: rdata <= W_Q3_0_0_3;
268: rdata <= W_Q3_0_0_4;
269: rdata <= W_Q3_0_0_5;
270: rdata <= W_Q3_0_0_6;
271: rdata <= W_Q3_0_0_7;
272: rdata <= W_Q3_0_1_0;
273: rdata <= W_Q3_0_1_1;
274: rdata <= W_Q3_0_1_2;
275: rdata <= W_Q3_0_1_3;
276: rdata <= W_Q3_0_1_4;
277: rdata <= W_Q3_0_1_5;
278: rdata <= W_Q3_0_1_6;
279: rdata <= W_Q3_0_1_7;
280: rdata <= W_Q3_1_0_0;
281: rdata <= W_Q3_1_0_1;
282: rdata <= W_Q3_1_0_2;
283: rdata <= W_Q3_1_0_3;
284: rdata <= W_Q3_1_1_0;
285: rdata <= W_Q3_1_1_1;
286: rdata <= W_Q3_1_1_2;
287: rdata <= W_Q3_1_1_3;
288: rdata <= W_Q3_1_2_0;
289: rdata <= W_Q3_1_2_1;
290: rdata <= W_Q3_1_2_2;
291: rdata <= W_Q3_1_2_3;
292: rdata <= W_Q3_1_3_0;
293: rdata <= W_Q3_1_3_1;
294: rdata <= W_Q3_1_3_2;
295: rdata <= W_Q3_1_3_3;
296: rdata <= W_Q3_1_4_0;
297: rdata <= W_Q3_1_4_1;
298: rdata <= W_Q3_1_4_2;
299: rdata <= W_Q3_1_4_3;
300: rdata <= W_Q3_1_5_0;
301: rdata <= W_Q3_1_5_1;
302: rdata <= W_Q3_1_5_2;
303: rdata <= W_Q3_1_5_3;
304: rdata <= W_Q3_1_6_0;
305: rdata <= W_Q3_1_6_1;
306: rdata <= W_Q3_1_6_2;
307: rdata <= W_Q3_1_6_3;
308: rdata <= W_Q3_1_7_0;
309: rdata <= W_Q3_1_7_1;
310: rdata <= W_Q3_1_7_2;
311: rdata <= W_Q3_1_7_3;
312: rdata <= W_Q3_2_0_0;
313: rdata <= W_Q3_2_1_0;
314: rdata <= W_Q3_2_2_0;
315: rdata <= W_Q3_2_3_0;
316: rdata <= B_Q3_0_0;
317: rdata <= B_Q3_0_1;
318: rdata <= B_Q3_0_2;
319: rdata <= B_Q3_0_3;
320: rdata <= B_Q3_0_4;
321: rdata <= B_Q3_0_5;
322: rdata <= B_Q3_0_6;
323: rdata <= B_Q3_0_7;
324: rdata <= B_Q3_1_0;
325: rdata <= B_Q3_1_1;
326: rdata <= B_Q3_1_2;
327: rdata <= B_Q3_1_3;
328: rdata <= B_Q3_2_0;
329: rdata <= W_Q4_0_0_0;
330: rdata <= W_Q4_0_0_1;
331: rdata <= W_Q4_0_0_2;
332: rdata <= W_Q4_0_0_3;
333: rdata <= W_Q4_0_0_4;
334: rdata <= W_Q4_0_0_5;
335: rdata <= W_Q4_0_0_6;
336: rdata <= W_Q4_0_0_7;
337: rdata <= W_Q4_0_1_0;
338: rdata <= W_Q4_0_1_1;
339: rdata <= W_Q4_0_1_2;
340: rdata <= W_Q4_0_1_3;
341: rdata <= W_Q4_0_1_4;
342: rdata <= W_Q4_0_1_5;
343: rdata <= W_Q4_0_1_6;
344: rdata <= W_Q4_0_1_7;
345: rdata <= W_Q4_1_0_0;
346: rdata <= W_Q4_1_0_1;
347: rdata <= W_Q4_1_0_2;
348: rdata <= W_Q4_1_0_3;
349: rdata <= W_Q4_1_1_0;
350: rdata <= W_Q4_1_1_1;
351: rdata <= W_Q4_1_1_2;
352: rdata <= W_Q4_1_1_3;
353: rdata <= W_Q4_1_2_0;
354: rdata <= W_Q4_1_2_1;
355: rdata <= W_Q4_1_2_2;
356: rdata <= W_Q4_1_2_3;
357: rdata <= W_Q4_1_3_0;
358: rdata <= W_Q4_1_3_1;
359: rdata <= W_Q4_1_3_2;
360: rdata <= W_Q4_1_3_3;
361: rdata <= W_Q4_1_4_0;
362: rdata <= W_Q4_1_4_1;
363: rdata <= W_Q4_1_4_2;
364: rdata <= W_Q4_1_4_3;
365: rdata <= W_Q4_1_5_0;
366: rdata <= W_Q4_1_5_1;
367: rdata <= W_Q4_1_5_2;
368: rdata <= W_Q4_1_5_3;
369: rdata <= W_Q4_1_6_0;
370: rdata <= W_Q4_1_6_1;
371: rdata <= W_Q4_1_6_2;
372: rdata <= W_Q4_1_6_3;
373: rdata <= W_Q4_1_7_0;
374: rdata <= W_Q4_1_7_1;
375: rdata <= W_Q4_1_7_2;
376: rdata <= W_Q4_1_7_3;
377: rdata <= W_Q4_2_0_0;
378: rdata <= W_Q4_2_1_0;
379: rdata <= W_Q4_2_2_0;
380: rdata <= W_Q4_2_3_0;
381: rdata <= B_Q4_0_0;
382: rdata <= B_Q4_0_1;
383: rdata <= B_Q4_0_2;
384: rdata <= B_Q4_0_3;
385: rdata <= B_Q4_0_4;
386: rdata <= B_Q4_0_5;
387: rdata <= B_Q4_0_6;
388: rdata <= B_Q4_0_7;
389: rdata <= B_Q4_1_0;
390: rdata <= B_Q4_1_1;
391: rdata <= B_Q4_1_2;
392: rdata <= B_Q4_1_3;
393: rdata <= B_Q4_2_0;
394: rdata <= W_Q5_0_0_0;
395: rdata <= W_Q5_0_0_1;
396: rdata <= W_Q5_0_0_2;
397: rdata <= W_Q5_0_0_3;
398: rdata <= W_Q5_0_0_4;
399: rdata <= W_Q5_0_0_5;
400: rdata <= W_Q5_0_0_6;
401: rdata <= W_Q5_0_0_7;
402: rdata <= W_Q5_0_1_0;
403: rdata <= W_Q5_0_1_1;
404: rdata <= W_Q5_0_1_2;
405: rdata <= W_Q5_0_1_3;
406: rdata <= W_Q5_0_1_4;
407: rdata <= W_Q5_0_1_5;
408: rdata <= W_Q5_0_1_6;
409: rdata <= W_Q5_0_1_7;
410: rdata <= W_Q5_1_0_0;
411: rdata <= W_Q5_1_0_1;
412: rdata <= W_Q5_1_0_2;
413: rdata <= W_Q5_1_0_3;
414: rdata <= W_Q5_1_1_0;
415: rdata <= W_Q5_1_1_1;
416: rdata <= W_Q5_1_1_2;
417: rdata <= W_Q5_1_1_3;
418: rdata <= W_Q5_1_2_0;
419: rdata <= W_Q5_1_2_1;
420: rdata <= W_Q5_1_2_2;
421: rdata <= W_Q5_1_2_3;
422: rdata <= W_Q5_1_3_0;
423: rdata <= W_Q5_1_3_1;
424: rdata <= W_Q5_1_3_2;
425: rdata <= W_Q5_1_3_3;
426: rdata <= W_Q5_1_4_0;
427: rdata <= W_Q5_1_4_1;
428: rdata <= W_Q5_1_4_2;
429: rdata <= W_Q5_1_4_3;
430: rdata <= W_Q5_1_5_0;
431: rdata <= W_Q5_1_5_1;
432: rdata <= W_Q5_1_5_2;
433: rdata <= W_Q5_1_5_3;
434: rdata <= W_Q5_1_6_0;
435: rdata <= W_Q5_1_6_1;
436: rdata <= W_Q5_1_6_2;
437: rdata <= W_Q5_1_6_3;
438: rdata <= W_Q5_1_7_0;
439: rdata <= W_Q5_1_7_1;
440: rdata <= W_Q5_1_7_2;
441: rdata <= W_Q5_1_7_3;
442: rdata <= W_Q5_2_0_0;
443: rdata <= W_Q5_2_1_0;
444: rdata <= W_Q5_2_2_0;
445: rdata <= W_Q5_2_3_0;
446: rdata <= B_Q5_0_0;
447: rdata <= B_Q5_0_1;
448: rdata <= B_Q5_0_2;
449: rdata <= B_Q5_0_3;
450: rdata <= B_Q5_0_4;
451: rdata <= B_Q5_0_5;
452: rdata <= B_Q5_0_6;
453: rdata <= B_Q5_0_7;
454: rdata <= B_Q5_1_0;
455: rdata <= B_Q5_1_1;
456: rdata <= B_Q5_1_2;
457: rdata <= B_Q5_1_3;
458: rdata <= B_Q5_2_0;
459: rdata <= W_Q6_0_0_0;
460: rdata <= W_Q6_0_0_1;
461: rdata <= W_Q6_0_0_2;
462: rdata <= W_Q6_0_0_3;
463: rdata <= W_Q6_0_0_4;
464: rdata <= W_Q6_0_0_5;
465: rdata <= W_Q6_0_0_6;
466: rdata <= W_Q6_0_0_7;
467: rdata <= W_Q6_0_1_0;
468: rdata <= W_Q6_0_1_1;
469: rdata <= W_Q6_0_1_2;
470: rdata <= W_Q6_0_1_3;
471: rdata <= W_Q6_0_1_4;
472: rdata <= W_Q6_0_1_5;
473: rdata <= W_Q6_0_1_6;
474: rdata <= W_Q6_0_1_7;
475: rdata <= W_Q6_1_0_0;
476: rdata <= W_Q6_1_0_1;
477: rdata <= W_Q6_1_0_2;
478: rdata <= W_Q6_1_0_3;
479: rdata <= W_Q6_1_1_0;
480: rdata <= W_Q6_1_1_1;
481: rdata <= W_Q6_1_1_2;
482: rdata <= W_Q6_1_1_3;
483: rdata <= W_Q6_1_2_0;
484: rdata <= W_Q6_1_2_1;
485: rdata <= W_Q6_1_2_2;
486: rdata <= W_Q6_1_2_3;
487: rdata <= W_Q6_1_3_0;
488: rdata <= W_Q6_1_3_1;
489: rdata <= W_Q6_1_3_2;
490: rdata <= W_Q6_1_3_3;
491: rdata <= W_Q6_1_4_0;
492: rdata <= W_Q6_1_4_1;
493: rdata <= W_Q6_1_4_2;
494: rdata <= W_Q6_1_4_3;
495: rdata <= W_Q6_1_5_0;
496: rdata <= W_Q6_1_5_1;
497: rdata <= W_Q6_1_5_2;
498: rdata <= W_Q6_1_5_3;
499: rdata <= W_Q6_1_6_0;
500: rdata <= W_Q6_1_6_1;
501: rdata <= W_Q6_1_6_2;
502: rdata <= W_Q6_1_6_3;
503: rdata <= W_Q6_1_7_0;
504: rdata <= W_Q6_1_7_1;
505: rdata <= W_Q6_1_7_2;
506: rdata <= W_Q6_1_7_3;
507: rdata <= W_Q6_2_0_0;
508: rdata <= W_Q6_2_1_0;
509: rdata <= W_Q6_2_2_0;
510: rdata <= W_Q6_2_3_0;
511: rdata <= B_Q6_0_0;
512: rdata <= B_Q6_0_1;
513: rdata <= B_Q6_0_2;
514: rdata <= B_Q6_0_3;
515: rdata <= B_Q6_0_4;
516: rdata <= B_Q6_0_5;
517: rdata <= B_Q6_0_6;
518: rdata <= B_Q6_0_7;
519: rdata <= B_Q6_1_0;
520: rdata <= B_Q6_1_1;
521: rdata <= B_Q6_1_2;
522: rdata <= B_Q6_1_3;
523: rdata <= B_Q6_2_0;
524: rdata <= W_Q7_0_0_0;
525: rdata <= W_Q7_0_0_1;
526: rdata <= W_Q7_0_0_2;
527: rdata <= W_Q7_0_0_3;
528: rdata <= W_Q7_0_0_4;
529: rdata <= W_Q7_0_0_5;
530: rdata <= W_Q7_0_0_6;
531: rdata <= W_Q7_0_0_7;
532: rdata <= W_Q7_0_1_0;
533: rdata <= W_Q7_0_1_1;
534: rdata <= W_Q7_0_1_2;
535: rdata <= W_Q7_0_1_3;
536: rdata <= W_Q7_0_1_4;
537: rdata <= W_Q7_0_1_5;
538: rdata <= W_Q7_0_1_6;
539: rdata <= W_Q7_0_1_7;
540: rdata <= W_Q7_1_0_0;
541: rdata <= W_Q7_1_0_1;
542: rdata <= W_Q7_1_0_2;
543: rdata <= W_Q7_1_0_3;
544: rdata <= W_Q7_1_1_0;
545: rdata <= W_Q7_1_1_1;
546: rdata <= W_Q7_1_1_2;
547: rdata <= W_Q7_1_1_3;
548: rdata <= W_Q7_1_2_0;
549: rdata <= W_Q7_1_2_1;
550: rdata <= W_Q7_1_2_2;
551: rdata <= W_Q7_1_2_3;
552: rdata <= W_Q7_1_3_0;
553: rdata <= W_Q7_1_3_1;
554: rdata <= W_Q7_1_3_2;
555: rdata <= W_Q7_1_3_3;
556: rdata <= W_Q7_1_4_0;
557: rdata <= W_Q7_1_4_1;
558: rdata <= W_Q7_1_4_2;
559: rdata <= W_Q7_1_4_3;
560: rdata <= W_Q7_1_5_0;
561: rdata <= W_Q7_1_5_1;
562: rdata <= W_Q7_1_5_2;
563: rdata <= W_Q7_1_5_3;
564: rdata <= W_Q7_1_6_0;
565: rdata <= W_Q7_1_6_1;
566: rdata <= W_Q7_1_6_2;
567: rdata <= W_Q7_1_6_3;
568: rdata <= W_Q7_1_7_0;
569: rdata <= W_Q7_1_7_1;
570: rdata <= W_Q7_1_7_2;
571: rdata <= W_Q7_1_7_3;
572: rdata <= W_Q7_2_0_0;
573: rdata <= W_Q7_2_1_0;
574: rdata <= W_Q7_2_2_0;
575: rdata <= W_Q7_2_3_0;
576: rdata <= B_Q7_0_0;
577: rdata <= B_Q7_0_1;
578: rdata <= B_Q7_0_2;
579: rdata <= B_Q7_0_3;
580: rdata <= B_Q7_0_4;
581: rdata <= B_Q7_0_5;
582: rdata <= B_Q7_0_6;
583: rdata <= B_Q7_0_7;
584: rdata <= B_Q7_1_0;
585: rdata <= B_Q7_1_1;
586: rdata <= B_Q7_1_2;
587: rdata <= B_Q7_1_3;
588: rdata <= B_Q7_2_0;
589: rdata <= min_Q0_I;
590: rdata <= min_Q0_Q;
591: rdata <= min_Q1_I;
592: rdata <= min_Q1_Q;
593: rdata <= min_Q2_I;
594: rdata <= min_Q2_Q;
595: rdata <= min_Q3_I;
596: rdata <= min_Q3_Q;
597: rdata <= min_Q4_I;
598: rdata <= min_Q4_Q;
599: rdata <= min_Q5_I;
600: rdata <= min_Q5_Q;
601: rdata <= min_Q6_I;
602: rdata <= min_Q6_Q;
603: rdata <= min_Q7_I;
604: rdata <= min_Q7_Q;
   default:rdata <= 32'hdeadbeef;
  endcase
 end
end
assign lb.rdata=rdata;
assign lb.rvalid=lb.rden16[READDELAY+1];
assign lb.rvalidlast=lb.rdenlast16[READDELAY+1];
endinterface