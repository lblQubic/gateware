	.aresetn( aresetn )
	,.pl_clk0( pl_clk0 )
,.cfgresetn00( cfgresetn00 )
,.cfgresetn01( cfgresetn01 )
,.cfgresetn02( cfgresetn02 )
,.cfgresetn03( cfgresetn03 )
,.cfgresetn04( cfgresetn04 )
,.cfgresetn05( cfgresetn05 )
,.cfgresetn06( cfgresetn06 )
,.cfgresetn07( cfgresetn07 )
,.cfgresetn08( cfgresetn08 )
,.cfgresetn09( cfgresetn09 )
,.cfgresetn10( cfgresetn10 )
,.cfgresetn11( cfgresetn11 )
,.cfgresetn12( cfgresetn12 )
,.cfgresetn13( cfgresetn13 )
,.cfgresetn14( cfgresetn14 )
,.cfgresetn15( cfgresetn15 )
,.cfgresetn16( cfgresetn16 )
,.cfgresetn17( cfgresetn17 )
,.cfgresetn18( cfgresetn18 )
,.dspresetn00( dspresetn00 )
,.dspresetn01( dspresetn01 )
,.dspresetn02( dspresetn02 )
,.dspresetn03( dspresetn03 )
,.dspresetn04( dspresetn04 )
,.dspresetn05( dspresetn05 )
,.dspresetn06( dspresetn06 )
,.dspresetn07( dspresetn07 )


,.psresetn00( psresetn00 )
,.psresetn01( psresetn01 )
,.psresetn02( psresetn02 )
,.adc2resetn00( adc2resetn00 )
,.adc2resetn01( adc2resetn01 )
,.adc2resetn02( adc2resetn02 )


,.lb1_wren( lb1_wren )
,.lb1_rden( lb1_rden )
,.lb1_waddr( lb1_waddr )
,.lb1_wdata( lb1_wdata )
,.lb1_raddr( lb1_raddr )
,.lb1_rdata( lb1_rdata )
,.lb1_rvalid( lb1_rvalid )
,.lb1_clk( lb1_clk )
,.lb1_aresetn( lb1_aresetn )
,.lb2_wren( lb2_wren )
,.lb2_rden( lb2_rden )
,.lb2_waddr( lb2_waddr )
,.lb2_wdata( lb2_wdata )
,.lb2_raddr( lb2_raddr )
,.lb2_rdata( lb2_rdata )
,.lb2_rvalid( lb2_rvalid )
,.lb2_clk( lb2_clk )
,.lb2_aresetn( lb2_aresetn )
,.BRAM_READ0_clk( BRAM_READ0_clk )
,.BRAM_READ0_rst( BRAM_READ0_rst )
,.BRAM_READ0_addr( BRAM_READ0_addr )
,.BRAM_READ0_din( BRAM_READ0_din )
,.BRAM_READ0_dout( BRAM_READ0_dout )
,.BRAM_READ0_en( BRAM_READ0_en )
,.BRAM_READ0_we( BRAM_READ0_we )
//,.bram_rsta_busy( bram_rsta_busy )
//,.bram_rstb_busy( bram_rstb_busy )
,.BRAM_READ1_clk( BRAM_READ1_clk )
,.BRAM_READ1_rst( BRAM_READ1_rst )
,.BRAM_READ1_addr( BRAM_READ1_addr )
,.BRAM_READ1_din( BRAM_READ1_din )
,.BRAM_READ1_dout( BRAM_READ1_dout )
,.BRAM_READ1_en( BRAM_READ1_en )
,.BRAM_READ1_we( BRAM_READ1_we )


,.BRAM_WRITE0_clk( BRAM_WRITE0_clk )
,.BRAM_WRITE0_rst( BRAM_WRITE0_rst )
,.BRAM_WRITE0_addr( BRAM_WRITE0_addr )
,.BRAM_WRITE0_din( BRAM_WRITE0_din )
,.BRAM_WRITE0_dout( BRAM_WRITE0_dout )
,.BRAM_WRITE0_en( BRAM_WRITE0_en )
,.BRAM_WRITE0_we( BRAM_WRITE0_we )
,.BRAM_WRITE1_clk( BRAM_WRITE1_clk )
,.BRAM_WRITE1_rst( BRAM_WRITE1_rst )
,.BRAM_WRITE1_addr( BRAM_WRITE1_addr )
,.BRAM_WRITE1_din( BRAM_WRITE1_din )
,.BRAM_WRITE1_dout( BRAM_WRITE1_dout )
,.BRAM_WRITE1_en( BRAM_WRITE1_en )
,.BRAM_WRITE1_we( BRAM_WRITE1_we )

,.BRAM_WRITE2_clk( BRAM_WRITE2_clk )
,.BRAM_WRITE2_rst( BRAM_WRITE2_rst )
,.BRAM_WRITE2_addr( BRAM_WRITE2_addr )
,.BRAM_WRITE2_din( BRAM_WRITE2_din )
,.BRAM_WRITE2_dout( BRAM_WRITE2_dout )
,.BRAM_WRITE2_en( BRAM_WRITE2_en )
,.BRAM_WRITE2_we( BRAM_WRITE2_we )
,.BRAM_WRITE3_clk( BRAM_WRITE3_clk )
,.BRAM_WRITE3_rst( BRAM_WRITE3_rst )
,.BRAM_WRITE3_addr( BRAM_WRITE3_addr )
,.BRAM_WRITE3_din( BRAM_WRITE3_din )
,.BRAM_WRITE3_dout( BRAM_WRITE3_dout )
,.BRAM_WRITE3_en( BRAM_WRITE3_en )
,.BRAM_WRITE3_we( BRAM_WRITE3_we )

,.clkadc2_300( clkadc2_300 )
,.clkadc2_600( clkadc2_600 )
,.DAC20_M_AXIS_ACLK( DAC20_M_AXIS_ACLK )
,.DAC20_M_AXIS_ARESETN( DAC20_M_AXIS_ARESETN )
,.DAC20_M_AXIS_TREADY( DAC20_M_AXIS_TREADY )
,.DAC20_M_AXIS_TVALID( DAC20_M_AXIS_TVALID )
,.DAC20_M_AXIS_TDATA( DAC20_M_AXIS_TDATA )
,.DAC20_M_AXIS_TSTRB( DAC20_M_AXIS_TSTRB )
,.DAC20_M_AXIS_TLAST( DAC20_M_AXIS_TLAST )
,.DAC22_M_AXIS_ACLK( DAC22_M_AXIS_ACLK )
,.DAC22_M_AXIS_ARESETN( DAC22_M_AXIS_ARESETN )
,.DAC22_M_AXIS_TREADY( DAC22_M_AXIS_TREADY )
,.DAC22_M_AXIS_TVALID( DAC22_M_AXIS_TVALID )
,.DAC22_M_AXIS_TDATA( DAC22_M_AXIS_TDATA )
,.DAC22_M_AXIS_TSTRB( DAC22_M_AXIS_TSTRB )
,.DAC22_M_AXIS_TLAST( DAC22_M_AXIS_TLAST )
,.clk_dac2( clk_dac2 )
,.DAC30_M_AXIS_ACLK( DAC30_M_AXIS_ACLK )
,.DAC30_M_AXIS_ARESETN( DAC30_M_AXIS_ARESETN )
,.DAC30_M_AXIS_TREADY( DAC30_M_AXIS_TREADY )
,.DAC30_M_AXIS_TVALID( DAC30_M_AXIS_TVALID )
,.DAC30_M_AXIS_TDATA( DAC30_M_AXIS_TDATA )
,.DAC30_M_AXIS_TSTRB( DAC30_M_AXIS_TSTRB )
,.DAC30_M_AXIS_TLAST( DAC30_M_AXIS_TLAST )
,.DAC32_M_AXIS_ACLK( DAC32_M_AXIS_ACLK )
,.DAC32_M_AXIS_ARESETN( DAC32_M_AXIS_ARESETN )
,.DAC32_M_AXIS_TREADY( DAC32_M_AXIS_TREADY )
,.DAC32_M_AXIS_TVALID( DAC32_M_AXIS_TVALID )
,.DAC32_M_AXIS_TDATA( DAC32_M_AXIS_TDATA )
,.DAC32_M_AXIS_TSTRB( DAC32_M_AXIS_TSTRB )
,.DAC32_M_AXIS_TLAST( DAC32_M_AXIS_TLAST )
,.clk_dac3( clk_dac3 )

,.ADC20_S_AXIS_ACLK( ADC20_S_AXIS_ACLK )
,.ADC20_S_AXIS_ARESETN( ADC20_S_AXIS_ARESETN )
,.ADC20_S_AXIS_TREADY( ADC20_S_AXIS_TREADY )
,.ADC20_S_AXIS_TVALID( ADC20_S_AXIS_TVALID )
,.ADC20_S_AXIS_TDATA( ADC20_S_AXIS_TDATA )
,.ADC20_S_AXIS_TSTRB( ADC20_S_AXIS_TSTRB )
,.ADC20_S_AXIS_TLAST( ADC20_S_AXIS_TLAST )
,.clk_adc2( clk_adc2 )
,.ADC21_S_AXIS_ACLK( ADC21_S_AXIS_ACLK )
,.ADC21_S_AXIS_ARESETN( ADC21_S_AXIS_ARESETN )
,.ADC21_S_AXIS_TREADY( ADC21_S_AXIS_TREADY )
,.ADC21_S_AXIS_TVALID( ADC21_S_AXIS_TVALID )
,.ADC21_S_AXIS_TDATA( ADC21_S_AXIS_TDATA )
,.ADC21_S_AXIS_TSTRB( ADC21_S_AXIS_TSTRB )
,.ADC21_S_AXIS_TLAST( ADC21_S_AXIS_TLAST )

,.cfgclk( cfgclk )
,.dspclk( dspclk )
