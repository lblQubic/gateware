output cfgresetn0
,output cfgresetn1
,output cfgresetn2
,output cfgresetn3
,output cfgresetn4
,output cfgresetn5
,output cfgresetn6
,output cfgresetn7
,output dspresetn0
,output dspresetn1
,output dspresetn2
,output dspresetn3
,output dspresetn4
,output dspresetn5
,output dspresetn6
,output dspresetn7
,output dspresetn8
,output dspresetn9
,output dspresetn10
,output dspresetn11
,output dspresetn12
,output dspresetn13
,output dspresetn14
,output dspresetn15
,output dspresetn16
,output dspresetn17
,output dspresetn18
,output dspresetn19
,output dspresetn20
,output dspresetn21
,output dspresetn22
,output dspresetn23
,output dspresetn24
,output dspresetn25
,output dspresetn26
,output dspresetn27
,output dspresetn28
,output dspresetn29
,output dspresetn30
,output dspresetn31
,output dspresetn32
,output dspresetn33
,output dspresetn34
,output dspresetn35
,output dspresetn36
,output dspresetn37
,output dspresetn38
,output dspresetn39
,output dspresetn40
,output dspresetn41
,output psresetn0
,output psresetn1
,output psresetn2
,output adc3resetn0