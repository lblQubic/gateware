interface ifdspregs #(parameter integer DATA_WIDTH = 32,parameter integer ADDR_WIDTH=24, parameter integer READDELAY=1)(    iflocalbus.lb lb
);
modport regs(input resetacc,stb_resetacc,amp,stb_amp,bramsel,stb_bramsel,coef00,stb_coef00,coef01,stb_coef01,coef02,stb_coef02,coef03,stb_coef03,coef10,stb_coef10,coef11,stb_coef11,coef12,stb_coef12,coef13,stb_coef13,coef20,stb_coef20,coef21,stb_coef21,coef22,stb_coef22,coef23,stb_coef23,coef30,stb_coef30,coef31,stb_coef31,coef32,stb_coef32,coef33,stb_coef33,dacsel,stb_dacsel,dspreset,stb_dspreset,nshot,stb_nshot,qdrvfreqsel,stb_qdrvfreqsel,rdlofreqsel,stb_rdlofreqsel,rdrvfreqsel,stb_rdrvfreqsel,reset_bram_read,stb_reset_bram_read,start,stb_start,test,stb_test,acqbufreset,stb_acqbufreset,dacmonreset,stb_dacmonreset,decimator,stb_decimator,acqchansel0,stb_acqchansel0,acqchansel1,stb_acqchansel1,dacmonchansel0,stb_dacmonchansel0,dacmonchansel1,stb_dacmonchansel1,dacmonchansel2,stb_dacmonchansel2,dacmonchansel3,stb_dacmonchansel3,delayaftertrig,stb_delayaftertrig,mixbb1sel,stb_mixbb1sel,mixbb2sel,stb_mixbb2sel,shift,stb_shift
,output addr_accbuf_mon0,addr_accbuf_mon1,addr_accbuf_mon2,addr_accbuf_mon3,busy,lastshotdone,shotcnt,test1,procdone,cnt00,cnt01,cnt02,cnt03,cnt10,cnt11,cnt12,cnt13,cnt20,cnt21,cnt22,cnt23,cnt30,cnt31,cnt32,cnt33
);
logic [DATA_WIDTH-1:0] rdata;
logic [DATA_WIDTH-1:0] wdata;
logic [ADDR_WIDTH-1:0] waddr;
logic [1-1:0] wren;

wire [32-1:0] resetacc;reg [32-1:0] reg_resetacc=0;reg stb_resetacc;assign resetacc=reg_resetacc;
wire [32-1:0] addr_accbuf_mon0;
wire [32-1:0] addr_accbuf_mon1;
wire [32-1:0] addr_accbuf_mon2;
wire [32-1:0] addr_accbuf_mon3;
wire [32-1:0] amp;reg [32-1:0] reg_amp=32000;reg stb_amp;assign amp=reg_amp;
wire [32-1:0] bramsel;reg [32-1:0] reg_bramsel=0;reg stb_bramsel;assign bramsel=reg_bramsel;
wire [4-1:0] busy;
wire [32-1:0] coef00;reg [32-1:0] reg_coef00=2147418112;reg stb_coef00;assign coef00=reg_coef00;
wire [32-1:0] coef01;reg [32-1:0] reg_coef01=0;reg stb_coef01;assign coef01=reg_coef01;
wire [32-1:0] coef02;reg [32-1:0] reg_coef02=0;reg stb_coef02;assign coef02=reg_coef02;
wire [32-1:0] coef03;reg [32-1:0] reg_coef03=0;reg stb_coef03;assign coef03=reg_coef03;
wire [32-1:0] coef10;reg [32-1:0] reg_coef10=0;reg stb_coef10;assign coef10=reg_coef10;
wire [32-1:0] coef11;reg [32-1:0] reg_coef11=2147418112;reg stb_coef11;assign coef11=reg_coef11;
wire [32-1:0] coef12;reg [32-1:0] reg_coef12=0;reg stb_coef12;assign coef12=reg_coef12;
wire [32-1:0] coef13;reg [32-1:0] reg_coef13=0;reg stb_coef13;assign coef13=reg_coef13;
wire [32-1:0] coef20;reg [32-1:0] reg_coef20=0;reg stb_coef20;assign coef20=reg_coef20;
wire [32-1:0] coef21;reg [32-1:0] reg_coef21=0;reg stb_coef21;assign coef21=reg_coef21;
wire [32-1:0] coef22;reg [32-1:0] reg_coef22=2147418112;reg stb_coef22;assign coef22=reg_coef22;
wire [32-1:0] coef23;reg [32-1:0] reg_coef23=0;reg stb_coef23;assign coef23=reg_coef23;
wire [32-1:0] coef30;reg [32-1:0] reg_coef30=0;reg stb_coef30;assign coef30=reg_coef30;
wire [32-1:0] coef31;reg [32-1:0] reg_coef31=0;reg stb_coef31;assign coef31=reg_coef31;
wire [32-1:0] coef32;reg [32-1:0] reg_coef32=0;reg stb_coef32;assign coef32=reg_coef32;
wire [32-1:0] coef33;reg [32-1:0] reg_coef33=2147418112;reg stb_coef33;assign coef33=reg_coef33;
wire [32-1:0] dacsel;reg [32-1:0] reg_dacsel=3;reg stb_dacsel;assign dacsel=reg_dacsel;
wire [1-1:0] dspreset;reg [1-1:0] reg_dspreset=0;reg stb_dspreset;assign dspreset=reg_dspreset;
wire [1-1:0] lastshotdone;
wire [32-1:0] nshot;reg [32-1:0] reg_nshot=10;reg stb_nshot;assign nshot=reg_nshot;
wire [32-1:0] qdrvfreqsel;reg [32-1:0] reg_qdrvfreqsel=3;reg stb_qdrvfreqsel;assign qdrvfreqsel=reg_qdrvfreqsel;
wire [32-1:0] rdlofreqsel;reg [32-1:0] reg_rdlofreqsel=3;reg stb_rdlofreqsel;assign rdlofreqsel=reg_rdlofreqsel;
wire [32-1:0] rdrvfreqsel;reg [32-1:0] reg_rdrvfreqsel=3;reg stb_rdrvfreqsel;assign rdrvfreqsel=reg_rdrvfreqsel;
wire [32-1:0] reset_bram_read;reg [32-1:0] reg_reset_bram_read=0;reg stb_reset_bram_read;assign reset_bram_read=reg_reset_bram_read;
wire [32-1:0] shotcnt;
wire [1-1:0] start;reg [1-1:0] reg_start=0;reg stb_start;assign start=reg_start;
wire [32-1:0] test;reg [32-1:0] reg_test=0;reg stb_test;assign test=reg_test;
wire [32-1:0] test1;
wire [1-1:0] acqbufreset;reg [1-1:0] reg_acqbufreset=1;reg stb_acqbufreset;assign acqbufreset=reg_acqbufreset;
wire [1-1:0] dacmonreset;reg [1-1:0] reg_dacmonreset=1;reg stb_dacmonreset;assign dacmonreset=reg_dacmonreset;
wire [8-1:0] decimator;reg [8-1:0] reg_decimator=1;reg stb_decimator;assign decimator=reg_decimator;
wire [5-1:0] acqchansel0;reg [5-1:0] reg_acqchansel0=1;reg stb_acqchansel0;assign acqchansel0=reg_acqchansel0;
wire [5-1:0] acqchansel1;reg [5-1:0] reg_acqchansel1=0;reg stb_acqchansel1;assign acqchansel1=reg_acqchansel1;
wire [5-1:0] dacmonchansel0;reg [5-1:0] reg_dacmonchansel0=0;reg stb_dacmonchansel0;assign dacmonchansel0=reg_dacmonchansel0;
wire [5-1:0] dacmonchansel1;reg [5-1:0] reg_dacmonchansel1=0;reg stb_dacmonchansel1;assign dacmonchansel1=reg_dacmonchansel1;
wire [5-1:0] dacmonchansel2;reg [5-1:0] reg_dacmonchansel2=0;reg stb_dacmonchansel2;assign dacmonchansel2=reg_dacmonchansel2;
wire [5-1:0] dacmonchansel3;reg [5-1:0] reg_dacmonchansel3=0;reg stb_dacmonchansel3;assign dacmonchansel3=reg_dacmonchansel3;
wire [16-1:0] delayaftertrig;reg [16-1:0] reg_delayaftertrig=100;reg stb_delayaftertrig;assign delayaftertrig=reg_delayaftertrig;
wire [16-1:0] mixbb1sel;reg [16-1:0] reg_mixbb1sel=0;reg stb_mixbb1sel;assign mixbb1sel=reg_mixbb1sel;
wire [16-1:0] mixbb2sel;reg [16-1:0] reg_mixbb2sel=1;reg stb_mixbb2sel;assign mixbb2sel=reg_mixbb2sel;
wire [5-1:0] shift;reg [5-1:0] reg_shift=15;reg stb_shift;assign shift=reg_shift;
wire [32-1:0] procdone;
wire [32-1:0] cnt00;
wire [32-1:0] cnt01;
wire [32-1:0] cnt02;
wire [32-1:0] cnt03;
wire [32-1:0] cnt10;
wire [32-1:0] cnt11;
wire [32-1:0] cnt12;
wire [32-1:0] cnt13;
wire [32-1:0] cnt20;
wire [32-1:0] cnt21;
wire [32-1:0] cnt22;
wire [32-1:0] cnt23;
wire [32-1:0] cnt30;
wire [32-1:0] cnt31;
wire [32-1:0] cnt32;
wire [32-1:0] cnt33;
always @(posedge lb.clk) begin
wdata<=lb.wdata;
waddr<=lb.waddr;
wren<=lb.wren;
stb_resetacc<=(lb.waddr==1)&lb.wren;if (stb_resetacc) reg_resetacc<=wdata[32-1:0];
stb_amp<=(lb.waddr==6)&lb.wren;if (stb_amp) reg_amp<=wdata[32-1:0];
stb_bramsel<=(lb.waddr==7)&lb.wren;if (stb_bramsel) reg_bramsel<=wdata[32-1:0];
stb_coef00<=(lb.waddr==9)&lb.wren;if (stb_coef00) reg_coef00<=wdata[32-1:0];
stb_coef01<=(lb.waddr==10)&lb.wren;if (stb_coef01) reg_coef01<=wdata[32-1:0];
stb_coef02<=(lb.waddr==11)&lb.wren;if (stb_coef02) reg_coef02<=wdata[32-1:0];
stb_coef03<=(lb.waddr==12)&lb.wren;if (stb_coef03) reg_coef03<=wdata[32-1:0];
stb_coef10<=(lb.waddr==13)&lb.wren;if (stb_coef10) reg_coef10<=wdata[32-1:0];
stb_coef11<=(lb.waddr==14)&lb.wren;if (stb_coef11) reg_coef11<=wdata[32-1:0];
stb_coef12<=(lb.waddr==15)&lb.wren;if (stb_coef12) reg_coef12<=wdata[32-1:0];
stb_coef13<=(lb.waddr==16)&lb.wren;if (stb_coef13) reg_coef13<=wdata[32-1:0];
stb_coef20<=(lb.waddr==17)&lb.wren;if (stb_coef20) reg_coef20<=wdata[32-1:0];
stb_coef21<=(lb.waddr==18)&lb.wren;if (stb_coef21) reg_coef21<=wdata[32-1:0];
stb_coef22<=(lb.waddr==19)&lb.wren;if (stb_coef22) reg_coef22<=wdata[32-1:0];
stb_coef23<=(lb.waddr==20)&lb.wren;if (stb_coef23) reg_coef23<=wdata[32-1:0];
stb_coef30<=(lb.waddr==21)&lb.wren;if (stb_coef30) reg_coef30<=wdata[32-1:0];
stb_coef31<=(lb.waddr==22)&lb.wren;if (stb_coef31) reg_coef31<=wdata[32-1:0];
stb_coef32<=(lb.waddr==23)&lb.wren;if (stb_coef32) reg_coef32<=wdata[32-1:0];
stb_coef33<=(lb.waddr==24)&lb.wren;if (stb_coef33) reg_coef33<=wdata[32-1:0];
stb_dacsel<=(lb.waddr==25)&lb.wren;if (stb_dacsel) reg_dacsel<=wdata[32-1:0];
stb_dspreset<=(lb.waddr==26)&lb.wren;if (stb_dspreset) reg_dspreset<=wdata[1-1:0];
stb_nshot<=(lb.waddr==28)&lb.wren;if (stb_nshot) reg_nshot<=wdata[32-1:0];
stb_qdrvfreqsel<=(lb.waddr==29)&lb.wren;if (stb_qdrvfreqsel) reg_qdrvfreqsel<=wdata[32-1:0];
stb_rdlofreqsel<=(lb.waddr==30)&lb.wren;if (stb_rdlofreqsel) reg_rdlofreqsel<=wdata[32-1:0];
stb_rdrvfreqsel<=(lb.waddr==31)&lb.wren;if (stb_rdrvfreqsel) reg_rdrvfreqsel<=wdata[32-1:0];
stb_reset_bram_read<=(lb.waddr==32)&lb.wren;if (stb_reset_bram_read) reg_reset_bram_read<=wdata[32-1:0];
stb_start<=(lb.waddr==34)&lb.wren;if (stb_start) reg_start<=wdata[1-1:0];
stb_test<=(lb.waddr==35)&lb.wren;if (stb_test) reg_test<=wdata[32-1:0];
stb_acqbufreset<=(lb.waddr==37)&lb.wren;if (stb_acqbufreset) reg_acqbufreset<=wdata[1-1:0];
stb_dacmonreset<=(lb.waddr==38)&lb.wren;if (stb_dacmonreset) reg_dacmonreset<=wdata[1-1:0];
stb_decimator<=(lb.waddr==39)&lb.wren;if (stb_decimator) reg_decimator<=wdata[8-1:0];
stb_acqchansel0<=(lb.waddr==40)&lb.wren;if (stb_acqchansel0) reg_acqchansel0<=wdata[5-1:0];
stb_acqchansel1<=(lb.waddr==41)&lb.wren;if (stb_acqchansel1) reg_acqchansel1<=wdata[5-1:0];
stb_dacmonchansel0<=(lb.waddr==42)&lb.wren;if (stb_dacmonchansel0) reg_dacmonchansel0<=wdata[5-1:0];
stb_dacmonchansel1<=(lb.waddr==43)&lb.wren;if (stb_dacmonchansel1) reg_dacmonchansel1<=wdata[5-1:0];
stb_dacmonchansel2<=(lb.waddr==44)&lb.wren;if (stb_dacmonchansel2) reg_dacmonchansel2<=wdata[5-1:0];
stb_dacmonchansel3<=(lb.waddr==45)&lb.wren;if (stb_dacmonchansel3) reg_dacmonchansel3<=wdata[5-1:0];
stb_delayaftertrig<=(lb.waddr==46)&lb.wren;if (stb_delayaftertrig) reg_delayaftertrig<=wdata[16-1:0];
stb_mixbb1sel<=(lb.waddr==47)&lb.wren;if (stb_mixbb1sel) reg_mixbb1sel<=wdata[16-1:0];
stb_mixbb2sel<=(lb.waddr==48)&lb.wren;if (stb_mixbb2sel) reg_mixbb2sel<=wdata[16-1:0];
stb_shift<=(lb.waddr==49)&lb.wren;if (stb_shift) reg_shift<=wdata[5-1:0];
end
always @(posedge lb.clk) begin
if (lb.rden16[READDELAY]) begin
case (lb.raddr16[(READDELAY+1)*ADDR_WIDTH-1:READDELAY*ADDR_WIDTH]) 

1: rdata <= resetacc;
2: rdata <= addr_accbuf_mon0;
3: rdata <= addr_accbuf_mon1;
4: rdata <= addr_accbuf_mon2;
5: rdata <= addr_accbuf_mon3;
6: rdata <= amp;
7: rdata <= bramsel;
8: rdata <= busy;
9: rdata <= coef00;
10: rdata <= coef01;
11: rdata <= coef02;
12: rdata <= coef03;
13: rdata <= coef10;
14: rdata <= coef11;
15: rdata <= coef12;
16: rdata <= coef13;
17: rdata <= coef20;
18: rdata <= coef21;
19: rdata <= coef22;
20: rdata <= coef23;
21: rdata <= coef30;
22: rdata <= coef31;
23: rdata <= coef32;
24: rdata <= coef33;
25: rdata <= dacsel;
26: rdata <= dspreset;
27: rdata <= lastshotdone;
28: rdata <= nshot;
29: rdata <= qdrvfreqsel;
30: rdata <= rdlofreqsel;
31: rdata <= rdrvfreqsel;
32: rdata <= reset_bram_read;
33: rdata <= shotcnt;
34: rdata <= start;
35: rdata <= test;
36: rdata <= test1;
37: rdata <= acqbufreset;
38: rdata <= dacmonreset;
39: rdata <= decimator;
40: rdata <= acqchansel0;
41: rdata <= acqchansel1;
42: rdata <= dacmonchansel0;
43: rdata <= dacmonchansel1;
44: rdata <= dacmonchansel2;
45: rdata <= dacmonchansel3;
46: rdata <= delayaftertrig;
47: rdata <= mixbb1sel;
48: rdata <= mixbb2sel;
49: rdata <= shift;
50: rdata <= procdone;
51: rdata <= cnt00;
52: rdata <= cnt01;
53: rdata <= cnt02;
54: rdata <= cnt03;
55: rdata <= cnt10;
56: rdata <= cnt11;
57: rdata <= cnt12;
58: rdata <= cnt13;
59: rdata <= cnt20;
60: rdata <= cnt21;
61: rdata <= cnt22;
62: rdata <= cnt23;
63: rdata <= cnt30;
64: rdata <= cnt31;
65: rdata <= cnt32;
66: rdata <= cnt33;
   default:rdata <= 32'hdeadbeef;
  endcase
 end
end
assign lb.rdata=rdata;
assign lb.rvalid=lb.rden16[READDELAY+1];
assign lb.rvalidlast=lb.rdenlast16[READDELAY+1];
endinterface