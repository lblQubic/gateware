module gitrevision(output [31:0] git);
assign git=32'h8ca7c80f;
endmodule
