.aresetn(aresetn)
,.pl_clk0(pl_clk0)
,`include "reset_portinst.vh"
,.lb1_wren(lb1_wren)
,.lb1_rden(lb1_rden)
,.lb1_rdenlast(lb1_rdenlast)
,.lb1_waddr(lb1_waddr)
,.lb1_wdata(lb1_wdata)
,.lb1_raddr(lb1_raddr)
,.lb1_rdata(lb1_rdata)
,.lb1_rvalid(lb1_rvalid)
,.lb1_rvalidlast(lb1_rvalidlast)
,.lb1_clk(lb1_clk)
,.lb1_aresetn(lb1_aresetn)
,.lb2_wren(lb2_wren)
,.lb2_rden(lb2_rden)
,.lb2_rdenlast(lb2_rdenlast)
,.lb2_waddr(lb2_waddr)
,.lb2_wdata(lb2_wdata)
,.lb2_raddr(lb2_raddr)
,.lb2_rdata(lb2_rdata)
,.lb2_rvalid(lb2_rvalid)
,.lb2_rvalidlast(lb2_rvalidlast)
,.lb2_clk(lb2_clk)
,.lb2_aresetn(lb2_aresetn)

,.lb3_wren(lb3_wren)
,.lb3_rden(lb3_rden)
,.lb3_rdenlast(lb3_rdenlast)
,.lb3_waddr(lb3_waddr)
,.lb3_wdata(lb3_wdata)
,.lb3_raddr(lb3_raddr)
,.lb3_rdata(lb3_rdata)
,.lb3_rvalid(lb3_rvalid)
,.lb3_rvalidlast(lb3_rvalidlast)
,.lb3_clk(lb3_clk)
,.lb3_aresetn(lb3_aresetn)


,.lb4_wren(lb4_wren)
,.lb4_rden(lb4_rden)
,.lb4_rdenlast(lb4_rdenlast)
,.lb4_waddr(lb4_waddr)
,.lb4_wdata(lb4_wdata)
,.lb4_raddr(lb4_raddr)
,.lb4_rdata(lb4_rdata)
,.lb4_rvalid(lb4_rvalid)
,.lb4_rvalidlast(lb4_rvalidlast)
,.lb4_clk(lb4_clk)
,.lb4_aresetn(lb4_aresetn)

,.clkadc3_300(clkadc3_300)
,.clkadc3_600(clkadc3_600)

,`include "rfdc_portinst.vh"
,.cfgclk(cfgclk)
,.dspclk(dspclk)
