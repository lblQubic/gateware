axi4stream.master dac00axis
,axi4stream.master dac01axis
,axi4stream.master dac02axis
,axi4stream.master dac03axis
,axi4stream.master dac10axis
,axi4stream.master dac11axis
,axi4stream.master dac12axis
,axi4stream.master dac13axis
,axi4stream.master dac20axis
,axi4stream.master dac21axis
,axi4stream.master dac22axis
,axi4stream.master dac23axis
,axi4stream.master dac30axis
,axi4stream.master dac31axis
,axi4stream.master dac32axis
,axi4stream.master dac33axis
,axi4stream.slave adc00axis
,axi4stream.slave adc01axis
,axi4stream.slave adc02axis
,axi4stream.slave adc03axis
,axi4stream.slave adc10axis
,axi4stream.slave adc11axis
,axi4stream.slave adc12axis
,axi4stream.slave adc13axis
,axi4stream.slave adc20axis
,axi4stream.slave adc21axis
,axi4stream.slave adc22axis
,axi4stream.slave adc23axis
,axi4stream.slave adc30axis
,axi4stream.slave adc31axis
,axi4stream.slave adc32axis
,axi4stream.slave adc33axis