parameter DEBUG="true"
,parameter integer LB_DATAWIDTH=32
,parameter integer LB_ADDRWIDTH=10
,parameter integer LB3_DATAWIDTH=32
,parameter integer LB3_ADDRWIDTH=20
,parameter integer DAC_AXIS_DATAWIDTH=256
,parameter integer ADC_AXIS_DATAWIDTH=64
,parameter integer BRAMADDRWIDTH=32
,`include "bram_para.vh"
