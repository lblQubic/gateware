.ACCBUF0_clk(ACCBUF0_clk)
,.ACCBUF0_rst(ACCBUF0_rst)
,.ACCBUF0_addr(ACCBUF0_addr)
,.ACCBUF0_din(ACCBUF0_din)
,.ACCBUF0_dout(ACCBUF0_dout)
,.ACCBUF0_en(ACCBUF0_en)
,.ACCBUF0_we(ACCBUF0_we)

,.ACCBUF1_clk(ACCBUF1_clk)
,.ACCBUF1_rst(ACCBUF1_rst)
,.ACCBUF1_addr(ACCBUF1_addr)
,.ACCBUF1_din(ACCBUF1_din)
,.ACCBUF1_dout(ACCBUF1_dout)
,.ACCBUF1_en(ACCBUF1_en)
,.ACCBUF1_we(ACCBUF1_we)

,.ACCBUF2_clk(ACCBUF2_clk)
,.ACCBUF2_rst(ACCBUF2_rst)
,.ACCBUF2_addr(ACCBUF2_addr)
,.ACCBUF2_din(ACCBUF2_din)
,.ACCBUF2_dout(ACCBUF2_dout)
,.ACCBUF2_en(ACCBUF2_en)
,.ACCBUF2_we(ACCBUF2_we)

,.ACQBUF0_clk(ACQBUF0_clk)
,.ACQBUF0_rst(ACQBUF0_rst)
,.ACQBUF0_addr(ACQBUF0_addr)
,.ACQBUF0_din(ACQBUF0_din)
,.ACQBUF0_dout(ACQBUF0_dout)
,.ACQBUF0_en(ACQBUF0_en)
,.ACQBUF0_we(ACQBUF0_we)

,.ACQBUF1_clk(ACQBUF1_clk)
,.ACQBUF1_rst(ACQBUF1_rst)
,.ACQBUF1_addr(ACQBUF1_addr)
,.ACQBUF1_din(ACQBUF1_din)
,.ACQBUF1_dout(ACQBUF1_dout)
,.ACQBUF1_en(ACQBUF1_en)
,.ACQBUF1_we(ACQBUF1_we)

,.COMMAND0_clk(COMMAND0_clk)
,.COMMAND0_rst(COMMAND0_rst)
,.COMMAND0_addr(COMMAND0_addr)
,.COMMAND0_din(COMMAND0_din)
,.COMMAND0_dout(COMMAND0_dout)
,.COMMAND0_en(COMMAND0_en)
,.COMMAND0_we(COMMAND0_we)

,.COMMAND1_clk(COMMAND1_clk)
,.COMMAND1_rst(COMMAND1_rst)
,.COMMAND1_addr(COMMAND1_addr)
,.COMMAND1_din(COMMAND1_din)
,.COMMAND1_dout(COMMAND1_dout)
,.COMMAND1_en(COMMAND1_en)
,.COMMAND1_we(COMMAND1_we)

,.COMMAND2_clk(COMMAND2_clk)
,.COMMAND2_rst(COMMAND2_rst)
,.COMMAND2_addr(COMMAND2_addr)
,.COMMAND2_din(COMMAND2_din)
,.COMMAND2_dout(COMMAND2_dout)
,.COMMAND2_en(COMMAND2_en)
,.COMMAND2_we(COMMAND2_we)

,.DACMON0_clk(DACMON0_clk)
,.DACMON0_rst(DACMON0_rst)
,.DACMON0_addr(DACMON0_addr)
,.DACMON0_din(DACMON0_din)
,.DACMON0_dout(DACMON0_dout)
,.DACMON0_en(DACMON0_en)
,.DACMON0_we(DACMON0_we)

,.DACMON1_clk(DACMON1_clk)
,.DACMON1_rst(DACMON1_rst)
,.DACMON1_addr(DACMON1_addr)
,.DACMON1_din(DACMON1_din)
,.DACMON1_dout(DACMON1_dout)
,.DACMON1_en(DACMON1_en)
,.DACMON1_we(DACMON1_we)

,.DACMON2_clk(DACMON2_clk)
,.DACMON2_rst(DACMON2_rst)
,.DACMON2_addr(DACMON2_addr)
,.DACMON2_din(DACMON2_din)
,.DACMON2_dout(DACMON2_dout)
,.DACMON2_en(DACMON2_en)
,.DACMON2_we(DACMON2_we)

,.DACMON3_clk(DACMON3_clk)
,.DACMON3_rst(DACMON3_rst)
,.DACMON3_addr(DACMON3_addr)
,.DACMON3_din(DACMON3_din)
,.DACMON3_dout(DACMON3_dout)
,.DACMON3_en(DACMON3_en)
,.DACMON3_we(DACMON3_we)

,.QDRVENV0_clk(QDRVENV0_clk)
,.QDRVENV0_rst(QDRVENV0_rst)
,.QDRVENV0_addr(QDRVENV0_addr)
,.QDRVENV0_din(QDRVENV0_din)
,.QDRVENV0_dout(QDRVENV0_dout)
,.QDRVENV0_en(QDRVENV0_en)
,.QDRVENV0_we(QDRVENV0_we)

,.QDRVENV1_clk(QDRVENV1_clk)
,.QDRVENV1_rst(QDRVENV1_rst)
,.QDRVENV1_addr(QDRVENV1_addr)
,.QDRVENV1_din(QDRVENV1_din)
,.QDRVENV1_dout(QDRVENV1_dout)
,.QDRVENV1_en(QDRVENV1_en)
,.QDRVENV1_we(QDRVENV1_we)

,.QDRVENV2_clk(QDRVENV2_clk)
,.QDRVENV2_rst(QDRVENV2_rst)
,.QDRVENV2_addr(QDRVENV2_addr)
,.QDRVENV2_din(QDRVENV2_din)
,.QDRVENV2_dout(QDRVENV2_dout)
,.QDRVENV2_en(QDRVENV2_en)
,.QDRVENV2_we(QDRVENV2_we)

,.QDRVFREQ0_clk(QDRVFREQ0_clk)
,.QDRVFREQ0_rst(QDRVFREQ0_rst)
,.QDRVFREQ0_addr(QDRVFREQ0_addr)
,.QDRVFREQ0_din(QDRVFREQ0_din)
,.QDRVFREQ0_dout(QDRVFREQ0_dout)
,.QDRVFREQ0_en(QDRVFREQ0_en)
,.QDRVFREQ0_we(QDRVFREQ0_we)

,.QDRVFREQ1_clk(QDRVFREQ1_clk)
,.QDRVFREQ1_rst(QDRVFREQ1_rst)
,.QDRVFREQ1_addr(QDRVFREQ1_addr)
,.QDRVFREQ1_din(QDRVFREQ1_din)
,.QDRVFREQ1_dout(QDRVFREQ1_dout)
,.QDRVFREQ1_en(QDRVFREQ1_en)
,.QDRVFREQ1_we(QDRVFREQ1_we)

,.QDRVFREQ2_clk(QDRVFREQ2_clk)
,.QDRVFREQ2_rst(QDRVFREQ2_rst)
,.QDRVFREQ2_addr(QDRVFREQ2_addr)
,.QDRVFREQ2_din(QDRVFREQ2_din)
,.QDRVFREQ2_dout(QDRVFREQ2_dout)
,.QDRVFREQ2_en(QDRVFREQ2_en)
,.QDRVFREQ2_we(QDRVFREQ2_we)

,.RDLOENV0_clk(RDLOENV0_clk)
,.RDLOENV0_rst(RDLOENV0_rst)
,.RDLOENV0_addr(RDLOENV0_addr)
,.RDLOENV0_din(RDLOENV0_din)
,.RDLOENV0_dout(RDLOENV0_dout)
,.RDLOENV0_en(RDLOENV0_en)
,.RDLOENV0_we(RDLOENV0_we)

,.RDLOENV1_clk(RDLOENV1_clk)
,.RDLOENV1_rst(RDLOENV1_rst)
,.RDLOENV1_addr(RDLOENV1_addr)
,.RDLOENV1_din(RDLOENV1_din)
,.RDLOENV1_dout(RDLOENV1_dout)
,.RDLOENV1_en(RDLOENV1_en)
,.RDLOENV1_we(RDLOENV1_we)

,.RDLOENV2_clk(RDLOENV2_clk)
,.RDLOENV2_rst(RDLOENV2_rst)
,.RDLOENV2_addr(RDLOENV2_addr)
,.RDLOENV2_din(RDLOENV2_din)
,.RDLOENV2_dout(RDLOENV2_dout)
,.RDLOENV2_en(RDLOENV2_en)
,.RDLOENV2_we(RDLOENV2_we)

,.RDLOFREQ0_clk(RDLOFREQ0_clk)
,.RDLOFREQ0_rst(RDLOFREQ0_rst)
,.RDLOFREQ0_addr(RDLOFREQ0_addr)
,.RDLOFREQ0_din(RDLOFREQ0_din)
,.RDLOFREQ0_dout(RDLOFREQ0_dout)
,.RDLOFREQ0_en(RDLOFREQ0_en)
,.RDLOFREQ0_we(RDLOFREQ0_we)

,.RDLOFREQ1_clk(RDLOFREQ1_clk)
,.RDLOFREQ1_rst(RDLOFREQ1_rst)
,.RDLOFREQ1_addr(RDLOFREQ1_addr)
,.RDLOFREQ1_din(RDLOFREQ1_din)
,.RDLOFREQ1_dout(RDLOFREQ1_dout)
,.RDLOFREQ1_en(RDLOFREQ1_en)
,.RDLOFREQ1_we(RDLOFREQ1_we)

,.RDLOFREQ2_clk(RDLOFREQ2_clk)
,.RDLOFREQ2_rst(RDLOFREQ2_rst)
,.RDLOFREQ2_addr(RDLOFREQ2_addr)
,.RDLOFREQ2_din(RDLOFREQ2_din)
,.RDLOFREQ2_dout(RDLOFREQ2_dout)
,.RDLOFREQ2_en(RDLOFREQ2_en)
,.RDLOFREQ2_we(RDLOFREQ2_we)

,.RDRVENV0_clk(RDRVENV0_clk)
,.RDRVENV0_rst(RDRVENV0_rst)
,.RDRVENV0_addr(RDRVENV0_addr)
,.RDRVENV0_din(RDRVENV0_din)
,.RDRVENV0_dout(RDRVENV0_dout)
,.RDRVENV0_en(RDRVENV0_en)
,.RDRVENV0_we(RDRVENV0_we)

,.RDRVENV1_clk(RDRVENV1_clk)
,.RDRVENV1_rst(RDRVENV1_rst)
,.RDRVENV1_addr(RDRVENV1_addr)
,.RDRVENV1_din(RDRVENV1_din)
,.RDRVENV1_dout(RDRVENV1_dout)
,.RDRVENV1_en(RDRVENV1_en)
,.RDRVENV1_we(RDRVENV1_we)

,.RDRVENV2_clk(RDRVENV2_clk)
,.RDRVENV2_rst(RDRVENV2_rst)
,.RDRVENV2_addr(RDRVENV2_addr)
,.RDRVENV2_din(RDRVENV2_din)
,.RDRVENV2_dout(RDRVENV2_dout)
,.RDRVENV2_en(RDRVENV2_en)
,.RDRVENV2_we(RDRVENV2_we)

,.RDRVFREQ0_clk(RDRVFREQ0_clk)
,.RDRVFREQ0_rst(RDRVFREQ0_rst)
,.RDRVFREQ0_addr(RDRVFREQ0_addr)
,.RDRVFREQ0_din(RDRVFREQ0_din)
,.RDRVFREQ0_dout(RDRVFREQ0_dout)
,.RDRVFREQ0_en(RDRVFREQ0_en)
,.RDRVFREQ0_we(RDRVFREQ0_we)

,.RDRVFREQ1_clk(RDRVFREQ1_clk)
,.RDRVFREQ1_rst(RDRVFREQ1_rst)
,.RDRVFREQ1_addr(RDRVFREQ1_addr)
,.RDRVFREQ1_din(RDRVFREQ1_din)
,.RDRVFREQ1_dout(RDRVFREQ1_dout)
,.RDRVFREQ1_en(RDRVFREQ1_en)
,.RDRVFREQ1_we(RDRVFREQ1_we)

,.RDRVFREQ2_clk(RDRVFREQ2_clk)
,.RDRVFREQ2_rst(RDRVFREQ2_rst)
,.RDRVFREQ2_addr(RDRVFREQ2_addr)
,.RDRVFREQ2_din(RDRVFREQ2_din)
,.RDRVFREQ2_dout(RDRVFREQ2_dout)
,.RDRVFREQ2_en(RDRVFREQ2_en)
,.RDRVFREQ2_we(RDRVFREQ2_we)
