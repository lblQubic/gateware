	.aresetn(aresetn)
	,.pl_clk0(pl_clk0)
,`include "reset_portinst.vh"
//,.cfgresetn00(cfgresetn00),.cfgresetn01(cfgresetn01),.cfgresetn02(cfgresetn02),.cfgresetn03(cfgresetn03),.cfgresetn04(cfgresetn04),.cfgresetn05(cfgresetn05),.cfgresetn06(cfgresetn06),.cfgresetn07(cfgresetn07)//,.cfgresetn08(cfgresetn08),.cfgresetn09(cfgresetn09)
//,.cfgresetn10(cfgresetn10),.cfgresetn11(cfgresetn11),.cfgresetn12(cfgresetn12),.cfgresetn13(cfgresetn13),.cfgresetn14(cfgresetn14),.cfgresetn15(cfgresetn15),.cfgresetn16(cfgresetn16),.cfgresetn17(cfgresetn17),.cfgresetn18(cfgresetn18),.cfgresetn19(cfgresetn19)
//,.cfgresetn20(cfgresetn20),.cfgresetn21(cfgresetn21),.cfgresetn22(cfgresetn22),.cfgresetn23(cfgresetn23),.cfgresetn24(cfgresetn24),.cfgresetn25(cfgresetn25),.cfgresetn26(cfgresetn26),.cfgresetn27(cfgresetn27),.cfgresetn28(cfgresetn28),.cfgresetn29(cfgresetn29)
//,.cfgresetn30(cfgresetn30),.cfgresetn31(cfgresetn31),.cfgresetn32(cfgresetn32),.cfgresetn33(cfgresetn33),.cfgresetn34(cfgresetn34),.cfgresetn35(cfgresetn35),.cfgresetn36(cfgresetn36),.cfgresetn37(cfgresetn37),.cfgresetn38(cfgresetn38),.cfgresetn39(cfgresetn39)
//,.cfgresetn40(cfgresetn40),.cfgresetn41(cfgresetn41),.cfgresetn42(cfgresetn42),.cfgresetn43(cfgresetn43),.cfgresetn44(cfgresetn44),.cfgresetn45(cfgresetn45),.cfgresetn46(cfgresetn46),.cfgresetn47(cfgresetn47),.cfgresetn48(cfgresetn48),.cfgresetn49(cfgresetn49)
//,.cfgresetn50(cfgresetn50),.cfgresetn51(cfgresetn51),.cfgresetn52(cfgresetn52),.cfgresetn53(cfgresetn53),.cfgresetn54(cfgresetn54),.cfgresetn55(cfgresetn55),.cfgresetn56(cfgresetn56),.cfgresetn57(cfgresetn57),.cfgresetn58(cfgresetn58),.cfgresetn59(cfgresetn59)
//,.cfgresetn60(cfgresetn60),.cfgresetn61(cfgresetn61),.cfgresetn62(cfgresetn62),.cfgresetn63(cfgresetn63),.cfgresetn64(cfgresetn64),.cfgresetn65(cfgresetn65),.cfgresetn66(cfgresetn66),.cfgresetn67(cfgresetn67),.cfgresetn68(cfgresetn68),.cfgresetn69(cfgresetn69)
//,.cfgresetn70(cfgresetn70),.cfgresetn71(cfgresetn71),.cfgresetn72(cfgresetn72),.cfgresetn73(cfgresetn73),.cfgresetn74(cfgresetn74),.cfgresetn75(cfgresetn75),.cfgresetn76(cfgresetn76),.cfgresetn77(cfgresetn77),.cfgresetn78(cfgresetn78),.cfgresetn79(cfgresetn79)
//,.cfgresetn80(cfgresetn80),.cfgresetn81(cfgresetn81),.cfgresetn82(cfgresetn82),.cfgresetn83(cfgresetn83),.cfgresetn84(cfgresetn84),.cfgresetn85(cfgresetn85),.cfgresetn86(cfgresetn86),.cfgresetn87(cfgresetn87),.cfgresetn88(cfgresetn88),.cfgresetn89(cfgresetn89)
//,.cfgresetn90(cfgresetn90),.cfgresetn91(cfgresetn91)

//,.dspresetn00(dspresetn00)
//,.dspresetn01(dspresetn01)
//,.dspresetn02(dspresetn02)
//,.dspresetn03(dspresetn03)
//,.dspresetn04(dspresetn04)
//,.dspresetn05(dspresetn05)
//,.dspresetn06(dspresetn06)
//,.dspresetn07(dspresetn07)
//
//
//,.psresetn00(psresetn00)
//,.psresetn01(psresetn01)
//,.psresetn02(psresetn02)
//,.adc2resetn00(adc2resetn00)
//,.adc2resetn01(adc2resetn01)
//,.adc2resetn02(adc2resetn02)
//

,.lb1_wren(lb1_wren)
,.lb1_rden(lb1_rden)
,.lb1_rdenlast(lb1_rdenlast)
,.lb1_waddr(lb1_waddr)
,.lb1_wdata(lb1_wdata)
,.lb1_raddr(lb1_raddr)
,.lb1_rdata(lb1_rdata)
,.lb1_rvalid(lb1_rvalid)
,.lb1_rvalidlast(lb1_rvalidlast)
,.lb1_clk(lb1_clk)
,.lb1_aresetn(lb1_aresetn)
,.lb2_wren(lb2_wren)
,.lb2_rden(lb2_rden)
,.lb2_rdenlast(lb2_rdenlast)
,.lb2_waddr(lb2_waddr)
,.lb2_wdata(lb2_wdata)
,.lb2_raddr(lb2_raddr)
,.lb2_rdata(lb2_rdata)
,.lb2_rvalid(lb2_rvalid)
,.lb2_rvalidlast(lb2_rvalidlast)
,.lb2_clk(lb2_clk)
,.lb2_aresetn(lb2_aresetn)

,.lb3_wren(lb3_wren)
,.lb3_rden(lb3_rden)
,.lb3_rdenlast(lb3_rdenlast)
,.lb3_waddr(lb3_waddr)
,.lb3_wdata(lb3_wdata)
,.lb3_raddr(lb3_raddr)
,.lb3_rdata(lb3_rdata)
,.lb3_rvalid(lb3_rvalid)
,.lb3_rvalidlast(lb3_rvalidlast)
,.lb3_clk(lb3_clk)
,.lb3_aresetn(lb3_aresetn)


,.lb4_wren(lb4_wren)
,.lb4_rden(lb4_rden)
,.lb4_rdenlast(lb4_rdenlast)
,.lb4_waddr(lb4_waddr)
,.lb4_wdata(lb4_wdata)
,.lb4_raddr(lb4_raddr)
,.lb4_rdata(lb4_rdata)
,.lb4_rvalid(lb4_rvalid)
,.lb4_rvalidlast(lb4_rvalidlast)
,.lb4_clk(lb4_clk)
,.lb4_aresetn(lb4_aresetn)

//,include "bram_portinst.vh"

,.clkadc2_300(clkadc2_300)
,.clkadc2_600(clkadc2_600)

/*,.DAC20_M_AXIS_ACLK(DAC20_M_AXIS_ACLK)
,.DAC20_M_AXIS_ARESETN(DAC20_M_AXIS_ARESETN)
,.DAC20_M_AXIS_TREADY(DAC20_M_AXIS_TREADY)
,.DAC20_M_AXIS_TVALID(DAC20_M_AXIS_TVALID)
,.DAC20_M_AXIS_TDATA(DAC20_M_AXIS_TDATA)
,.DAC20_M_AXIS_TSTRB(DAC20_M_AXIS_TSTRB)
,.DAC20_M_AXIS_TLAST(DAC20_M_AXIS_TLAST)
,.DAC22_M_AXIS_ACLK(DAC22_M_AXIS_ACLK)
,.DAC22_M_AXIS_ARESETN(DAC22_M_AXIS_ARESETN)
,.DAC22_M_AXIS_TREADY(DAC22_M_AXIS_TREADY)
,.DAC22_M_AXIS_TVALID(DAC22_M_AXIS_TVALID)
,.DAC22_M_AXIS_TDATA(DAC22_M_AXIS_TDATA)
,.DAC22_M_AXIS_TSTRB(DAC22_M_AXIS_TSTRB)
,.DAC22_M_AXIS_TLAST(DAC22_M_AXIS_TLAST)
,.clk_dac2(clk_dac2)
,.DAC30_M_AXIS_ACLK(DAC30_M_AXIS_ACLK)
,.DAC30_M_AXIS_ARESETN(DAC30_M_AXIS_ARESETN)
,.DAC30_M_AXIS_TREADY(DAC30_M_AXIS_TREADY)
,.DAC30_M_AXIS_TVALID(DAC30_M_AXIS_TVALID)
,.DAC30_M_AXIS_TDATA(DAC30_M_AXIS_TDATA)
,.DAC30_M_AXIS_TSTRB(DAC30_M_AXIS_TSTRB)
,.DAC30_M_AXIS_TLAST(DAC30_M_AXIS_TLAST)
,.DAC32_M_AXIS_ACLK(DAC32_M_AXIS_ACLK)
,.DAC32_M_AXIS_ARESETN(DAC32_M_AXIS_ARESETN)
,.DAC32_M_AXIS_TREADY(DAC32_M_AXIS_TREADY)
,.DAC32_M_AXIS_TVALID(DAC32_M_AXIS_TVALID)
,.DAC32_M_AXIS_TDATA(DAC32_M_AXIS_TDATA)
,.DAC32_M_AXIS_TSTRB(DAC32_M_AXIS_TSTRB)
,.DAC32_M_AXIS_TLAST(DAC32_M_AXIS_TLAST)
,.clk_dac3(clk_dac3)

,.ADC20_S_AXIS_ACLK(ADC20_S_AXIS_ACLK)
,.ADC20_S_AXIS_ARESETN(ADC20_S_AXIS_ARESETN)
,.ADC20_S_AXIS_TREADY(ADC20_S_AXIS_TREADY)
,.ADC20_S_AXIS_TVALID(ADC20_S_AXIS_TVALID)
,.ADC20_S_AXIS_TDATA(ADC20_S_AXIS_TDATA)
,.ADC20_S_AXIS_TSTRB(ADC20_S_AXIS_TSTRB)
,.ADC20_S_AXIS_TLAST(ADC20_S_AXIS_TLAST)
,.clk_adc2(clk_adc2)
,.ADC21_S_AXIS_ACLK(ADC21_S_AXIS_ACLK)
,.ADC21_S_AXIS_ARESETN(ADC21_S_AXIS_ARESETN)
,.ADC21_S_AXIS_TREADY(ADC21_S_AXIS_TREADY)
,.ADC21_S_AXIS_TVALID(ADC21_S_AXIS_TVALID)
,.ADC21_S_AXIS_TDATA(ADC21_S_AXIS_TDATA)
,.ADC21_S_AXIS_TSTRB(ADC21_S_AXIS_TSTRB)
,.ADC21_S_AXIS_TLAST(ADC21_S_AXIS_TLAST)
*/
,`include "rfdc_portinst.vh"
,.cfgclk(cfgclk)
,.dspclk(dspclk)
