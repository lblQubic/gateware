parameter integer ACCBUF_R_ADDRWIDTH=11,parameter integer ACCBUF_R_DATAWIDTH=32,parameter integer ACCBUF_R_DEPTH=2048,parameter integer ACCBUF_W_ADDRWIDTH=10,parameter integer ACCBUF_W_DATAWIDTH=64,parameter integer ACCBUF_W_DEPTH=1024
,parameter integer ACQBUF_R_ADDRWIDTH=13,parameter integer ACQBUF_R_DATAWIDTH=32,parameter integer ACQBUF_R_DEPTH=8192,parameter integer ACQBUF_W_ADDRWIDTH=12,parameter integer ACQBUF_W_DATAWIDTH=64,parameter integer ACQBUF_W_DEPTH=4096
,parameter integer COMMAND_R_ADDRWIDTH=11,parameter integer COMMAND_R_DATAWIDTH=128,parameter integer COMMAND_R_DEPTH=2048,parameter integer COMMAND_W_ADDRWIDTH=13,parameter integer COMMAND_W_DATAWIDTH=32,parameter integer COMMAND_W_DEPTH=8192
,parameter integer DACMON_R_ADDRWIDTH=12,parameter integer DACMON_R_DATAWIDTH=32,parameter integer DACMON_R_DEPTH=4096,parameter integer DACMON_W_ADDRWIDTH=9,parameter integer DACMON_W_DATAWIDTH=256,parameter integer DACMON_W_DEPTH=512
,parameter integer QDRVENV_R_ADDRWIDTH=8,parameter integer QDRVENV_R_DATAWIDTH=512,parameter integer QDRVENV_R_DEPTH=256,parameter integer QDRVENV_W_ADDRWIDTH=12,parameter integer QDRVENV_W_DATAWIDTH=32,parameter integer QDRVENV_W_DEPTH=4096
,parameter integer QDRVFREQ_R_ADDRWIDTH=9,parameter integer QDRVFREQ_R_DATAWIDTH=512,parameter integer QDRVFREQ_R_DEPTH=512,parameter integer QDRVFREQ_W_ADDRWIDTH=13,parameter integer QDRVFREQ_W_DATAWIDTH=32,parameter integer QDRVFREQ_W_DEPTH=8192
,parameter integer RDLOENV_R_ADDRWIDTH=12,parameter integer RDLOENV_R_DATAWIDTH=32,parameter integer RDLOENV_R_DEPTH=4096,parameter integer RDLOENV_W_ADDRWIDTH=12,parameter integer RDLOENV_W_DATAWIDTH=32,parameter integer RDLOENV_W_DEPTH=4096
,parameter integer RDLOFREQ_R_ADDRWIDTH=9,parameter integer RDLOFREQ_R_DATAWIDTH=128,parameter integer RDLOFREQ_R_DEPTH=512,parameter integer RDLOFREQ_W_ADDRWIDTH=11,parameter integer RDLOFREQ_W_DATAWIDTH=32,parameter integer RDLOFREQ_W_DEPTH=2048
,parameter integer RDRVENV_R_ADDRWIDTH=12,parameter integer RDRVENV_R_DATAWIDTH=32,parameter integer RDRVENV_R_DEPTH=4096,parameter integer RDRVENV_W_ADDRWIDTH=12,parameter integer RDRVENV_W_DATAWIDTH=32,parameter integer RDRVENV_W_DEPTH=4096
,parameter integer RDRVFREQ_R_ADDRWIDTH=9,parameter integer RDRVFREQ_R_DATAWIDTH=512,parameter integer RDRVFREQ_R_DEPTH=512,parameter integer RDRVFREQ_W_ADDRWIDTH=13,parameter integer RDRVFREQ_W_DATAWIDTH=32,parameter integer RDRVFREQ_W_DEPTH=8192
,parameter integer SDBUF_R_ADDRWIDTH=10,parameter integer SDBUF_R_DATAWIDTH=32,parameter integer SDBUF_R_DEPTH=1024,parameter integer SDBUF_W_ADDRWIDTH=10,parameter integer SDBUF_W_DATAWIDTH=32,parameter integer SDBUF_W_DEPTH=1024
,parameter integer SDPARA_R_ADDRWIDTH=7,parameter integer SDPARA_R_DATAWIDTH=32,parameter integer SDPARA_R_DEPTH=128,parameter integer SDPARA_W_ADDRWIDTH=7,parameter integer SDPARA_W_DATAWIDTH=32,parameter integer SDPARA_W_DEPTH=128