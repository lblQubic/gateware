ifbram acqbuf0_R
,ifbram acqbuf1_R
,ifbram command0_W
,ifbram command1_W
,ifbram command2_W
,ifbram command3_W
,ifbram command4_W
,ifbram command5_W
,ifbram command6_W
,ifbram command7_W
,ifbram qdrvfreq0_W
,ifbram qdrvfreq1_W
,ifbram qdrvfreq2_W
,ifbram qdrvfreq3_W
,ifbram qdrvfreq4_W
,ifbram qdrvfreq5_W
,ifbram qdrvfreq6_W
,ifbram qdrvfreq7_W
,ifbram rdrvfreq0_W
,ifbram rdrvfreq1_W
,ifbram rdrvfreq2_W
,ifbram rdrvfreq3_W
,ifbram rdrvfreq4_W
,ifbram rdrvfreq5_W
,ifbram rdrvfreq6_W
,ifbram rdrvfreq7_W
,ifbram dacmon0_R
,ifbram dacmon1_R
,ifbram dacmon2_R
,ifbram dacmon3_R
,ifbram qdrvenv0_W
,ifbram qdrvenv1_W
,ifbram qdrvenv2_W
,ifbram qdrvenv3_W
,ifbram qdrvenv4_W
,ifbram qdrvenv5_W
,ifbram qdrvenv6_W
,ifbram qdrvenv7_W
,ifbram rdloenv0_W
,ifbram rdloenv1_W
,ifbram rdloenv2_W
,ifbram rdloenv3_W
,ifbram rdloenv4_W
,ifbram rdloenv5_W
,ifbram rdloenv6_W
,ifbram rdloenv7_W
,ifbram rdrvenv0_W
,ifbram rdrvenv1_W
,ifbram rdrvenv2_W
,ifbram rdrvenv3_W
,ifbram rdrvenv4_W
,ifbram rdrvenv5_W
,ifbram rdrvenv6_W
,ifbram rdrvenv7_W
,ifbram accbuf0_R
,ifbram accbuf1_R
,ifbram accbuf2_R
,ifbram accbuf3_R
,ifbram accbuf4_R
,ifbram accbuf5_R
,ifbram accbuf6_R
,ifbram accbuf7_R
,ifbram rdlofreq0_W
,ifbram rdlofreq1_W
,ifbram rdlofreq2_W
,ifbram rdlofreq3_W
,ifbram rdlofreq4_W
,ifbram rdlofreq5_W
,ifbram rdlofreq6_W
,ifbram rdlofreq7_W
,ifbram sdbuf0_R
,ifbram sdbuf1_R
,ifbram sdbuf2_R
,ifbram sdbuf3_R
,ifbram sdbuf4_R
,ifbram sdbuf5_R
,ifbram sdbuf6_R
,ifbram sdbuf7_R
,ifbram sdpara0_W
,ifbram sdpara1_W
,ifbram sdpara2_W
,ifbram sdpara3_W
,ifbram sdpara4_W
,ifbram sdpara5_W
,ifbram sdpara6_W
,ifbram sdpara7_W