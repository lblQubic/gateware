localparam INITLMKADC={{4'h0,8'h2,8'h20,8'h0}
,{4'h0,8'h2,8'h0,8'h0}
,{4'h0,8'h2,8'h20,8'h0}
,{4'h2,8'h2,16'h2082}
,{4'h0,8'h3,8'h0,8'h0}
,{4'h0,8'h3,8'h6,8'h0}
,{4'h0,8'h3,8'h8,8'h0}
,{4'h0,8'h1,8'hf0,8'h0}
,{4'h0,8'h3,8'h0,8'h0}
,{4'h0,8'h3,8'h1,8'h0}
,{4'h0,8'h3,8'h8,8'h0}
,{4'h0,8'h1,8'hf0,8'h0}
,{4'h1,16'h0,8'h90}
,{4'h1,16'h0,8'h10}
,{4'h1,16'h0,8'h10}
,{4'h1,16'h148,8'h33}
,{4'h1,16'h0,8'h90}
,{4'h1,16'h0,8'h10}
,{4'h1,16'h0,8'h10}
,{4'h1,16'h100,8'h61}
,{4'h1,16'h101,8'h22}
,{4'h1,16'h103,8'h2}
,{4'h1,16'h104,8'h20}
,{4'h1,16'h106,8'hf0}
,{4'h1,16'h107,8'h55}
,{4'h1,16'h108,8'h64}
,{4'h1,16'h109,8'h22}
,{4'h1,16'h10b,8'h5}
,{4'h1,16'h10c,8'h20}
,{4'h1,16'h10e,8'hb0}
,{4'h1,16'h10f,8'h11}
,{4'h1,16'h110,8'h61}
,{4'h1,16'h111,8'h22}
,{4'h1,16'h113,8'h2}
,{4'h1,16'h114,8'h20}
,{4'h1,16'h116,8'hf0}
,{4'h1,16'h117,8'h57}
,{4'h1,16'h118,8'h61}
,{4'h1,16'h119,8'h22}
,{4'h1,16'h11b,8'h2}
,{4'h1,16'h11c,8'h20}
,{4'h1,16'h11e,8'hf0}
,{4'h1,16'h11f,8'h57}
,{4'h1,16'h120,8'h62}
,{4'h1,16'h121,8'h22}
,{4'h1,16'h123,8'h5}
,{4'h1,16'h124,8'h20}
,{4'h1,16'h126,8'hb0}
,{4'h1,16'h127,8'h11}
,{4'h1,16'h128,8'h68}
,{4'h1,16'h129,8'h22}
,{4'h1,16'h12c,8'h20}
,{4'h1,16'h12e,8'hf7}
,{4'h1,16'h12f,8'h1}
,{4'h1,16'h130,8'h61}
,{4'h1,16'h133,8'h2}
,{4'h1,16'h134,8'h20}
,{4'h1,16'h136,8'hf7}
,{4'h1,16'h138,8'h40}
,{4'h1,16'h139,8'h5}
,{4'h1,16'h13e,8'h0}
,{4'h1,16'h140,8'hf7}
,{4'h1,16'h143,8'h10}
,{4'h1,16'h144,8'hff}
,{4'h1,16'h145,8'h7f}
,{4'h1,16'h147,8'h10}
,{4'h1,16'h148,8'h33}
,{4'h1,16'h149,8'h0}
,{4'h1,16'h14a,8'h0}
,{4'h1,16'h14b,8'h5}
,{4'h1,16'h14c,8'hff}
,{4'h1,16'h150,8'h0}
,{4'h1,16'h156,8'h78}
,{4'h1,16'h15f,8'hb}
,{4'h1,16'h161,8'h1}
,{4'h1,16'h162,8'h44}
,{4'h1,16'h16e,8'h13}
,{4'h1,16'h173,8'h60}
,{4'h1,16'h1ffd,8'h0}
,{4'h1,16'h1ffe,8'h0}
,{4'h1,16'h1fff,8'h53}
,{4'h3,16'h11,8'h80}
,{4'h4,16'h11,8'h80}
,{4'h3,16'h53,8'h20}
,{4'h4,16'h53,8'h20}
,{4'h3,16'h59,8'h20}
,{4'h4,16'h59,8'h20}
,{4'h3,16'h4005,8'h0}
,{4'h4,16'h4005,8'h0}
,{4'h3,16'h4003,8'h0}
,{4'h4,16'h4003,8'h0}
,{4'h3,16'h4004,8'h69}
,{4'h4,16'h4004,8'h69}
,{4'h3,16'h6000,8'h80}
,{4'h4,16'h6000,8'h80}
,{4'h3,16'h6001,8'h4}
,{4'h4,16'h6001,8'h4}
,{4'h3,16'h6002,8'h0}
,{4'h4,16'h6002,8'h0}
,{4'h3,16'h6007,8'h8}
,{4'h4,16'h6007,8'h8}
,{4'h3,16'h4003,8'h0}
,{4'h4,16'h4003,8'h0}
,{4'h3,16'h4004,8'h6a}
,{4'h4,16'h4004,8'h6a}
,{4'h3,16'h6016,8'h2}
,{4'h4,16'h6016,8'h2}
,{4'h3,16'h6017,8'h40}
,{4'h4,16'h6017,8'h40}
,{4'h3,16'h6017,8'h0}
,{4'h4,16'h6017,8'h0}
,{4'h3,16'h4003,8'h0}
,{4'h4,16'h4003,8'h0}
,{4'h3,16'h4004,8'h68}
,{4'h4,16'h4004,8'h68}
,{4'h3,16'h6000,8'h1}
,{4'h4,16'h6000,8'h1}
,{4'h3,16'h6000,8'h0}
,{4'h4,16'h6000,8'h0}
,{4'h3,16'h4003,8'h0}
,{4'h4,16'h4003,8'h0}
,{4'h3,16'h4004,8'h69}
,{4'h4,16'h4004,8'h69}
,{4'h3,16'h6006,8'h1f}
,{4'h4,16'h6006,8'h1f}
,{4'h8,8'h2,8'h20,8'h0}
,{4'h8,8'h2,8'h0,8'h0}
,{4'h8,8'h2,8'h20,8'h0}
,{4'ha,8'h2,16'h2082}
,{4'h8,8'h3,8'h0,8'h0}
,{4'h8,8'h3,8'h6,8'h0}
,{4'h8,8'h3,8'h8,8'h0}
,{4'h8,8'h1,8'hf0,8'h0}
,{4'h8,8'h3,8'h0,8'h0}
,{4'h8,8'h3,8'h1,8'h0}
,{4'h8,8'h3,8'h8,8'h0}
,{4'h8,8'h1,8'hf0,8'h0}
,{4'h9,16'h0,8'h90}
,{4'h9,16'h0,8'h10}
,{4'h9,16'h0,8'h10}
,{4'h9,16'h148,8'h33}
,{4'h9,16'h0,8'h90}
,{4'h9,16'h0,8'h10}
,{4'h9,16'h0,8'h10}
,{4'h9,16'h100,8'h61}
,{4'h9,16'h101,8'h22}
,{4'h9,16'h103,8'h2}
,{4'h9,16'h104,8'h20}
,{4'h9,16'h106,8'hf0}
,{4'h9,16'h107,8'h55}
,{4'h9,16'h108,8'h64}
,{4'h9,16'h109,8'h22}
,{4'h9,16'h10b,8'h5}
,{4'h9,16'h10c,8'h20}
,{4'h9,16'h10e,8'hb0}
,{4'h9,16'h10f,8'h11}
,{4'h9,16'h110,8'h61}
,{4'h9,16'h111,8'h22}
,{4'h9,16'h113,8'h2}
,{4'h9,16'h114,8'h20}
,{4'h9,16'h116,8'hf0}
,{4'h9,16'h117,8'h57}
,{4'h9,16'h118,8'h61}
,{4'h9,16'h119,8'h22}
,{4'h9,16'h11b,8'h2}
,{4'h9,16'h11c,8'h20}
,{4'h9,16'h11e,8'hf0}
,{4'h9,16'h11f,8'h57}
,{4'h9,16'h120,8'h62}
,{4'h9,16'h121,8'h22}
,{4'h9,16'h123,8'h5}
,{4'h9,16'h124,8'h20}
,{4'h9,16'h126,8'hb0}
,{4'h9,16'h127,8'h11}
,{4'h9,16'h128,8'h68}
,{4'h9,16'h129,8'h22}
,{4'h9,16'h12c,8'h20}
,{4'h9,16'h12e,8'hf7}
,{4'h9,16'h12f,8'h1}
,{4'h9,16'h130,8'h61}
,{4'h9,16'h133,8'h2}
,{4'h9,16'h134,8'h20}
,{4'h9,16'h136,8'hf7}
,{4'h9,16'h138,8'h40}
,{4'h9,16'h139,8'h5}
,{4'h9,16'h13e,8'h0}
,{4'h9,16'h140,8'hf7}
,{4'h9,16'h143,8'h10}
,{4'h9,16'h144,8'hff}
,{4'h9,16'h145,8'h7f}
,{4'h9,16'h147,8'h10}
,{4'h9,16'h148,8'h33}
,{4'h9,16'h149,8'h0}
,{4'h9,16'h14a,8'h0}
,{4'h9,16'h14b,8'h5}
,{4'h9,16'h14c,8'hff}
,{4'h9,16'h150,8'h0}
,{4'h9,16'h156,8'h78}
,{4'h9,16'h15f,8'hb}
,{4'h9,16'h161,8'h1}
,{4'h9,16'h162,8'h44}
,{4'h9,16'h16e,8'h13}
,{4'h9,16'h173,8'h60}
,{4'h9,16'h1ffd,8'h0}
,{4'h9,16'h1ffe,8'h0}
,{4'h9,16'h1fff,8'h53}
,{4'hb,16'h11,8'h80}
,{4'hc,16'h11,8'h80}
,{4'hb,16'h53,8'h20}
,{4'hc,16'h53,8'h20}
,{4'hb,16'h59,8'h20}
,{4'hc,16'h59,8'h20}
,{4'hb,16'h4005,8'h0}
,{4'hc,16'h4005,8'h0}
,{4'hb,16'h4003,8'h0}
,{4'hc,16'h4003,8'h0}
,{4'hb,16'h4004,8'h69}
,{4'hc,16'h4004,8'h69}
,{4'hb,16'h6000,8'h80}
,{4'hc,16'h6000,8'h80}
,{4'hb,16'h6001,8'h4}
,{4'hc,16'h6001,8'h4}
,{4'hb,16'h6002,8'h0}
,{4'hc,16'h6002,8'h0}
,{4'hb,16'h6007,8'h8}
,{4'hc,16'h6007,8'h8}
,{4'hb,16'h4003,8'h0}
,{4'hc,16'h4003,8'h0}
,{4'hb,16'h4004,8'h6a}
,{4'hc,16'h4004,8'h6a}
,{4'hb,16'h6016,8'h2}
,{4'hc,16'h6016,8'h2}
,{4'hb,16'h6017,8'h40}
,{4'hc,16'h6017,8'h40}
,{4'hb,16'h6017,8'h0}
,{4'hc,16'h6017,8'h0}
,{4'hb,16'h4003,8'h0}
,{4'hc,16'h4003,8'h0}
,{4'hb,16'h4004,8'h68}
,{4'hc,16'h4004,8'h68}
,{4'hb,16'h6000,8'h1}
,{4'hc,16'h6000,8'h1}
,{4'hb,16'h6000,8'h0}
,{4'hc,16'h6000,8'h0}
,{4'hb,16'h4003,8'h0}
,{4'hc,16'h4003,8'h0}
,{4'hb,16'h4004,8'h69}
,{4'hc,16'h4004,8'h69}
,{4'hb,16'h6006,8'h1f}
,{4'hc,16'h6006,8'h1f}};
localparam INITDAC={{4'h2,8'h0,16'h18}
,{4'h2,8'h4a,16'hff1e}
,{4'h2,8'h1,16'ha0}
,{4'h2,8'h2,16'h2082}
,{4'h2,8'h1a,16'h20}
,{4'h2,8'h1e,16'h4444}
,{4'h2,8'h1f,16'h4440}
,{4'h2,8'h20,16'h4044}
,{4'h2,8'h24,16'h20}
,{4'h2,8'h25,16'h2000}
,{4'h2,8'h3b,16'h800}
,{4'h2,8'h3c,16'h228}
,{4'h2,8'h3e,16'h108}
,{4'h2,8'h4b,16'h0}
,{4'h2,8'h4c,16'h1f07}
,{4'h2,8'h4d,16'h300}
,{4'h2,8'h4e,16'hf4f}
,{4'h2,8'h51,16'hdf}
,{4'h2,8'h61,16'h1}
,{4'h2,8'h4a,16'hff1f}
,{4'h2,8'h4a,16'hff01}
,{4'ha,8'h0,16'h18}
,{4'ha,8'h4a,16'hff1e}
,{4'ha,8'h1,16'ha0}
,{4'ha,8'h2,16'h2082}
,{4'ha,8'h1a,16'h20}
,{4'ha,8'h1e,16'h4444}
,{4'ha,8'h1f,16'h4440}
,{4'ha,8'h20,16'h4044}
,{4'ha,8'h24,16'h20}
,{4'ha,8'h25,16'h2000}
,{4'ha,8'h3b,16'h800}
,{4'ha,8'h3c,16'h228}
,{4'ha,8'h3e,16'h108}
,{4'ha,8'h4b,16'h0}
,{4'ha,8'h4c,16'h1f07}
,{4'ha,8'h4d,16'h300}
,{4'ha,8'h4e,16'hf4f}
,{4'ha,8'h51,16'hdf}
,{4'ha,8'h61,16'h1}
,{4'ha,8'h4a,16'hff1f}
,{4'ha,8'h4a,16'hff01}};
localparam INITDAC2={
{4'h2,8'h4a,16'hff1f}
,{4'h2,8'h4a,16'hff01}
,{4'ha,8'h4a,16'hff1f}
,{4'ha,8'h4a,16'hff01}
};
localparam INITDAC2LEN=4;
localparam INITLMKADCLEN=250;
localparam INITDACLEN=42;
localparam I2CINITCMD= {{1'h1,4'h2,32'he8080000}
,{1'h0,4'h2,32'ha8000000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8010000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8020000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8030000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8040000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8050000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8060000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8070000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8080000}
,{1'h1,4'h2,32'ha9000000}
,{1'h0,4'h2,32'ha8090000}
,{1'h1,4'h2,32'ha9000000}
,{1'h1,4'h2,32'he8010000}
,{1'h1,4'h3,32'hba891000}
,{1'h1,4'h3,32'hba070300}
,{1'h1,4'h3,32'hba084300}
,{1'h1,4'h3,32'hba091000}
,{1'h1,4'h3,32'hba0a0100}
,{1'h1,4'h3,32'hba0bbd00}
,{1'h1,4'h3,32'hba0cf200}
,{1'h1,4'h3,32'hba890000}
,{1'h1,4'h3,32'hba874000}
,{1'h1,4'h2,32'he8800000}
,{1'h1,4'h3,32'hd0001400}
,{1'h1,4'h3,32'hd001e400}
,{1'h1,4'h3,32'hd002a200}
,{1'h1,4'h3,32'hd0031500}
,{1'h1,4'h3,32'hd0049200}
,{1'h1,4'h3,32'hd005ed00}
,{1'h1,4'h3,32'hd0062d00}
,{1'h1,4'h3,32'hd0072a00}
,{1'h1,4'h3,32'hd0080000}
,{1'h1,4'h3,32'hd009c000}
,{1'h1,4'h3,32'hd00a0800}
,{1'h1,4'h3,32'hd00b4200}
,{1'h1,4'h3,32'hd0132900}
,{1'h1,4'h3,32'hd0143e00}
,{1'h1,4'h3,32'hd015ff00}
,{1'h1,4'h3,32'hd016df00}
,{1'h1,4'h3,32'hd0171f00}
,{1'h1,4'h3,32'hd0183f00}
,{1'h1,4'h3,32'hd0192000}
,{1'h1,4'h3,32'hd01f0000}
,{1'h1,4'h3,32'hd0200000}
,{1'h1,4'h3,32'hd0210700}
,{1'h1,4'h3,32'hd0220000}
,{1'h1,4'h3,32'hd0230000}
,{1'h1,4'h3,32'hd0240700}
,{1'h1,4'h3,32'hd0286000}
,{1'h1,4'h3,32'hd0290100}
,{1'h1,4'h3,32'hd02a6700}
,{1'h1,4'h3,32'hd02b0000}
,{1'h1,4'h3,32'hd02c0000}
,{1'h1,4'h3,32'hd02d3e00}
,{1'h1,4'h3,32'hd02e0000}
,{1'h1,4'h3,32'hd02f0000}
,{1'h1,4'h3,32'hd0303e00}
,{1'h1,4'h3,32'hd0370000}
,{1'h1,4'h3,32'hd0831f00}
,{1'h1,4'h3,32'hd0840200}
,{1'h1,4'h3,32'hd0890100}
,{1'h1,4'h3,32'hd08a0f00}
,{1'h1,4'h3,32'hd08bff00}
,{1'h1,4'h3,32'hd08e0000}
,{1'h1,4'h3,32'hd08f0000}
,{1'h1,4'h3,32'hd0884000}
};
localparam I2CCMDLENGTH=75;

localparam AXIINITCMDLENGTH=20;
localparam AXIINITCMD={
{3'h0,12'h10,32'h101}
,{3'h0,12'h30,32'h1}
,{3'h0,12'h34,32'h1}
,{3'h1,12'h10,32'h101}
,{3'h1,12'h30,32'h1}
,{3'h1,12'h34,32'h1}
,{3'h2,12'h10,32'h101}
,{3'h2,12'h34,32'h1}
,{3'h2,12'h810,32'hf0f03}
,{3'h2,12'h814,32'h80000000}
,{3'h3,12'h10,32'h101}
,{3'h3,12'h30,32'h1}
,{3'h3,12'h34,32'h1}
,{3'h4,12'h10,32'h101}
,{3'h4,12'h30,32'h1}
,{3'h4,12'h34,32'h1}
,{3'h5,12'h10,32'h101}
,{3'h5,12'h34,32'h1}
,{3'h5,12'h810,32'hf0f03}
,{3'h5,12'h814,32'h80000000}
};
