module gteth_gt #(parameter GT_SIM_GTRESET_SPEEDUP = "TRUE",
parameter RX_DFE_KL_CFG2_IN = 32'h301148AC,
parameter PMA_RSV_IN = 32'h00018480,
parameter PCS_RSVD_ATTR_IN = 48'h000000000000
)(
output GTXTXN
,output GTXTXP
,input GTXRXP
,input GTXRXN
,input GTNORTHREFCLK0
,input GTNORTHREFCLK1
,input GTREFCLK0
,input GTREFCLK1
,input GTSOUTHREFCLK0
,input GTSOUTHREFCLK1
,input QPLLCLK
,input QPLLREFCLK
,input CPLLLOCKDETCLK
,input [2:0] CPLLREFCLKSEL


,input RXUSERRDY
,input TXUSERRDY
,input [15:0] TXDATA
,input [1:0] TXCHARISK
,output RXVALID
,output [15:0] RXDATA
,output [1:0] RXCHARISK
,output txusrclk
,output rxusrclk
,output txusrclk2
,output rxusrclk2
,input reset
,input readyforreset
,output resetdone
);
wire [47:0] rxdata_dummy;
wire [5:0] rxchariscomma_float_i;
wire [5:0] rxcharisk_float_i;
wire [5:0] rxdisperr_float_i;
wire [5:0] rxnotintable_float_i;
//wire resetalign;
wire txrxreset1;
wire txrxreset0;
wire txrxreset=txrxreset0|txrxreset1;
wire txcharisk=~resetdone ? 8'h1 : {6'h0,TXCHARISK};
wire [63:0] txdata=~resetdone ? 64'h000000bc : {32'b0,TXDATA} ;
wire CPLLRESET;
wire GTTXRESET=txrxreset;
wire GTRXRESET=txrxreset;
wire RXPMARESET=txrxreset;
wire RXRESETDONE;
wire TXRESETDONE;
wire [1:0] RXDISPERR;
wire [1:0] RXNOTINTABLE;
wire [1:0] RXCHARISCOMMA;
assign dbrxcharisk=RXCHARISK;
wire RXBYTEISALIGNED;
wire RXBYTEREALIGN;
wire RXCOMMADET;
wire CPLLLOCK;
wire CPLLFBCLKLOST;
wire CPLLREFCLKLOST;
wire RXOUTCLK;
wire TXUSRCLK;
wire TXUSRCLK2;
wire TXOUTCLK;
wire RXUSRCLK;
wire RXUSRCLK2;

GTXE2_CHANNEL #(.SIM_RECEIVER_DETECT_PASS("TRUE"),.SIM_TX_EIDLE_DRIVE_LEVEL("X"),.SIM_RESET_SPEEDUP(GT_SIM_GTRESET_SPEEDUP),.SIM_CPLLREFCLK_SEL(3'b001),.SIM_VERSION("4.0"),.ALIGN_COMMA_DOUBLE("FALSE"),.ALIGN_COMMA_ENABLE(10'b0001111111),.ALIGN_COMMA_WORD(2),.ALIGN_MCOMMA_DET("TRUE"),.ALIGN_MCOMMA_VALUE(10'b1010000011),.ALIGN_PCOMMA_DET("TRUE"),.ALIGN_PCOMMA_VALUE(10'b0101111100),.SHOW_REALIGN_COMMA("TRUE"),.RXSLIDE_AUTO_WAIT(7),.RXSLIDE_MODE("OFF"),.RX_SIG_VALID_DLY(10),.RX_DISPERR_SEQ_MATCH("TRUE"),.DEC_MCOMMA_DETECT("TRUE"),.DEC_PCOMMA_DETECT("TRUE"),.DEC_VALID_COMMA_ONLY("FALSE"),.CBCC_DATA_SOURCE_SEL("DECODED"),.CLK_COR_SEQ_2_USE("FALSE"),.CLK_COR_KEEP_IDLE("FALSE"),.CLK_COR_MAX_LAT(36),.CLK_COR_MIN_LAT(32),.CLK_COR_PRECEDENCE("TRUE"),.CLK_COR_REPEAT_WAIT(0),.CLK_COR_SEQ_LEN(1),.CLK_COR_SEQ_1_ENABLE(4'b1111),.CLK_COR_SEQ_1_1(10'b0100000000),.CLK_COR_SEQ_1_2(10'b0000000000),.CLK_COR_SEQ_1_3(10'b0000000000),.CLK_COR_SEQ_1_4(10'b0000000000),.CLK_CORRECT_USE("FALSE"),.CLK_COR_SEQ_2_ENABLE(4'b1111),.CLK_COR_SEQ_2_1(10'b0100000000),.CLK_COR_SEQ_2_2(10'b0000000000),.CLK_COR_SEQ_2_3(10'b0000000000),.CLK_COR_SEQ_2_4(10'b0000000000),.CHAN_BOND_KEEP_ALIGN("FALSE"),.CHAN_BOND_MAX_SKEW(1),.CHAN_BOND_SEQ_LEN(1),.CHAN_BOND_SEQ_1_1(10'b0000000000),.CHAN_BOND_SEQ_1_2(10'b0000000000),.CHAN_BOND_SEQ_1_3(10'b0000000000),.CHAN_BOND_SEQ_1_4(10'b0000000000),.CHAN_BOND_SEQ_1_ENABLE(4'b1111),.CHAN_BOND_SEQ_2_1(10'b0000000000),.CHAN_BOND_SEQ_2_2(10'b0000000000),.CHAN_BOND_SEQ_2_3(10'b0000000000),.CHAN_BOND_SEQ_2_4(10'b0000000000),.CHAN_BOND_SEQ_2_ENABLE(4'b1111),.CHAN_BOND_SEQ_2_USE("FALSE"),.FTS_DESKEW_SEQ_ENABLE(4'b1111),.FTS_LANE_DESKEW_CFG(4'b1111),.FTS_LANE_DESKEW_EN("FALSE"),.ES_CONTROL(6'b000000),.ES_ERRDET_EN("FALSE"),.ES_EYE_SCAN_EN("TRUE"),.ES_HORZ_OFFSET(12'h000),.ES_PMA_CFG(10'b0000000000),.ES_PRESCALE(5'b00000),.ES_QUALIFIER(80'h00000000000000000000),.ES_QUAL_MASK(80'h00000000000000000000),.ES_SDATA_MASK(80'h00000000000000000000),.ES_VERT_OFFSET(9'b000000000),.RX_DATA_WIDTH(20),.OUTREFCLK_SEL_INV(2'b11),.PMA_RSV(PMA_RSV_IN),.PMA_RSV2(16'h2050),.PMA_RSV3(2'b00),.PMA_RSV4(32'h00000000),.RX_BIAS_CFG(12'b000000000100),.DMONITOR_CFG(24'h000A00),.RX_CM_SEL(2'b11),.RX_CM_TRIM(3'b010),.RX_DEBUG_CFG(12'b000000000000),.RX_OS_CFG(13'b0000010000000),.TERM_RCAL_CFG(5'b10000),.TERM_RCAL_OVRD(1'b0),.TST_RSV(32'h00000000),.RX_CLK25_DIV(5),.TX_CLK25_DIV(5),.UCODEER_CLR(1'b0),.PCS_PCIE_EN("FALSE"),.PCS_RSVD_ATTR(PCS_RSVD_ATTR_IN),.RXBUF_ADDR_MODE("FAST"),.RXBUF_EIDLE_HI_CNT(4'b1000),.RXBUF_EIDLE_LO_CNT(4'b0000),.RXBUF_EN("TRUE"),.RX_BUFFER_CFG(6'b000000),.RXBUF_RESET_ON_CB_CHANGE("TRUE"),.RXBUF_RESET_ON_COMMAALIGN("FALSE"),.RXBUF_RESET_ON_EIDLE("FALSE"),.RXBUF_RESET_ON_RATE_CHANGE("TRUE"),.RXBUFRESET_TIME(5'b00001),.RXBUF_THRESH_OVFLW(61),.RXBUF_THRESH_OVRD("FALSE"),.RXBUF_THRESH_UNDFLW(8),.RXDLY_CFG(16'h001F),.RXDLY_LCFG(9'h030),.RXDLY_TAP_CFG(16'h0000),.RXPH_CFG(24'h000000),.RXPHDLY_CFG(24'h084020),.RXPH_MONITOR_SEL(5'b00000),.RX_XCLK_SEL("RXREC"),.RX_DDI_SEL(6'b000000),.RX_DEFER_RESET_BUF_EN("TRUE"),.RXCDR_CFG(72'h03000023ff10100020),.CPLL_FBDIV(4),.RXOUT_DIV(4),.TXOUT_DIV(4),.RXCDR_FR_RESET_ON_EIDLE(1'b0),.RXCDR_HOLD_DURING_EIDLE(1'b0),.RXCDR_PH_RESET_ON_EIDLE(1'b0),.RXCDR_LOCK_CFG(6'b010101),.RXCDRFREQRESET_TIME(5'b00001),.RXCDRPHRESET_TIME(5'b00001),.RXISCANRESET_TIME(5'b00001),.RXPCSRESET_TIME(5'b00001),.RXPMARESET_TIME(5'b00011),.RXOOB_CFG(7'b0000110),.RXGEARBOX_EN("FALSE"),.GEARBOX_MODE(3'b000),.RXPRBS_ERR_LOOPBACK(1'b0),.PD_TRANS_TIME_FROM_P2(12'h03c),.PD_TRANS_TIME_NONE_P2(8'h19),.PD_TRANS_TIME_TO_P2(8'h64),.SAS_MAX_COM(64),.SAS_MIN_COM(36),.SATA_BURST_SEQ_LEN(4'b0101),.SATA_BURST_VAL(3'b100),.SATA_EIDLE_VAL(3'b100),.SATA_MAX_BURST(8),.SATA_MAX_INIT(21),.SATA_MAX_WAKE(7),.SATA_MIN_BURST(4),.SATA_MIN_INIT(12),.SATA_MIN_WAKE(4),.TRANS_TIME_RATE(8'h0E),.TXBUF_EN("TRUE"),.TXBUF_RESET_ON_RATE_CHANGE("TRUE"),.TXDLY_CFG(16'h001F),.TXDLY_LCFG(9'h030),.TXDLY_TAP_CFG(16'h0000),.TXPH_CFG(16'h0780),.TXPHDLY_CFG(24'h084020),.TXPH_MONITOR_SEL(5'b00000),.TX_XCLK_SEL("TXOUT"),.TX_DATA_WIDTH(20),.TX_DEEMPH0(5'b00000),.TX_DEEMPH1(5'b00000),.TX_EIDLE_ASSERT_DELAY(3'b110),.TX_EIDLE_DEASSERT_DELAY(3'b100),.TX_LOOPBACK_DRIVE_HIZ("FALSE"),.TX_MAINCURSOR_SEL(1'b0),.TX_DRIVE_MODE("DIRECT"),.TX_MARGIN_FULL_0(7'b1001110),.TX_MARGIN_FULL_1(7'b1001001),.TX_MARGIN_FULL_2(7'b1000101),.TX_MARGIN_FULL_3(7'b1000010),.TX_MARGIN_FULL_4(7'b1000000),.TX_MARGIN_LOW_0(7'b1000110),.TX_MARGIN_LOW_1(7'b1000100),.TX_MARGIN_LOW_2(7'b1000010),.TX_MARGIN_LOW_3(7'b1000000),.TX_MARGIN_LOW_4(7'b1000000),.TXGEARBOX_EN("FALSE"),.TXPCSRESET_TIME(5'b00001),.TXPMARESET_TIME(5'b00001),.TX_RXDETECT_CFG(14'h1832),.TX_RXDETECT_REF(3'b100),.CPLL_CFG(24'hBC07DC),.CPLL_FBDIV_45(5),.CPLL_INIT_CFG(24'h00001E),.CPLL_LOCK_CFG(16'h01E8),.CPLL_REFCLK_DIV(1),.SATA_CPLL_CFG("VCO_3000MHZ"),.RXDFELPMRESET_TIME(7'b0001111),.RXLPM_HF_CFG(14'b00000011110000),.RXLPM_LF_CFG(14'b00000011110000),.RX_DFE_GAIN_CFG(23'h020FEA),.RX_DFE_H2_CFG(12'b000000000000),.RX_DFE_H3_CFG(12'b000001000000),.RX_DFE_H4_CFG(11'b00011110000),.RX_DFE_H5_CFG(11'b00011100000),.RX_DFE_KL_CFG(13'b0000011111110),.RX_DFE_LPM_CFG(16'h0904),.RX_DFE_LPM_HOLD_DURING_EIDLE(1'b0),.RX_DFE_UT_CFG(17'b10001111000000000),.RX_DFE_VP_CFG(17'b00011111100000011),.RX_CLKMUX_PD(1'b1),.TX_CLKMUX_PD(1'b1),.RX_INT_DATAWIDTH(0),.TX_INT_DATAWIDTH(0),.TX_QPI_STATUS_EN(1'b0),.RX_DFE_KL_CFG2(RX_DFE_KL_CFG2_IN),.RX_DFE_XYD_CFG(13'b0000000000000),.TX_PREDRIVER_MODE(1'b0))
GTXE2_CHANNEL(.CPLLLOCKEN(1'b1),.GTRSVD(16'b0000000000000000),.PCSRSVDIN(16'b0000000000000000),.PCSRSVDIN2(5'b00000),.PMARSVDIN(5'b00000),.PMARSVDIN2(5'b00000),.TSTIN(20'b11111111111111111111),.TSTOUT(),.CLKRSVD(4'b0),.GTGREFCLK(1'b0),.DRPADDR(9'b0),.DRPCLK(1'b0),.DRPDI(16'b0),.DRPDO(),.DRPEN(1'b0),.DRPRDY(),.DRPWE(1'b0),.GTREFCLKMONITOR(),.RXSYSCLKSEL(2'b00),.TXSYSCLKSEL(2'b00),.DMONITOROUT(),.TX8B10BEN(1'b1),.LOOPBACK(3'b0),.PHYSTATUS(),.RXRATE(3'b0),.RXPD(2'b0),.TXPD(2'b0),.SETERRSTATUS(1'b0),.EYESCANRESET(1'b0),.EYESCANDATAERROR(),.EYESCANMODE(1'b0),.EYESCANTRIGGER(),.RXCDRFREQRESET(1'b0),.RXCDRHOLD(1'b0),.RXCDRLOCK(),.RXCDROVRDEN(1'b0),.RXCDRRESET(1'b0),.RXCDRRESETRSV(1'b0),.RXCLKCORCNT(),.RX8B10BEN(1'b1),.RXPRBSERR(),.RXPRBSSEL(3'b0),.RXPRBSCNTRESET(1'b0),.RXDFEXYDEN(1'b1),.RXDFEXYDHOLD(1'b0),.RXDFEXYDOVRDEN(1'b0),.RXBUFRESET(1'b0),.RXBUFSTATUS(),.RXDDIEN(1'b0),.RXDLYBYPASS(1'b1),.RXDLYEN(1'b0),.RXDLYOVRDEN(1'b0),.RXDLYSRESET(1'b0),.RXDLYSRESETDONE(),.RXPHALIGN(1'b0),.RXPHALIGNDONE(),.RXPHALIGNEN(1'b0),.RXPHDLYPD(1'b0),.RXPHDLYRESET(1'b0),.RXPHMONITOR(),.RXPHOVRDEN(1'b0),.RXPHSLIPMONITOR(),.RXSTATUS(),.RXCOMMADETEN(1'b1),.RXCHANBONDSEQ(),.RXCHBONDEN(1'b0),.RXCHBONDLEVEL(3'b0),.RXCHBONDMASTER(1'b0),.RXCHBONDO(),.RXCHBONDSLAVE(1'b0),.RXCHANISALIGNED(),.RXCHANREALIGN(),.RXLPMHFHOLD(1'b0),.RXLPMHFOVRDEN(1'b0),.RXLPMLFHOLD(1'b0),.RXDFEAGCHOLD(1'b0),.RXDFEAGCOVRDEN(1'b0),.RXDFECM1EN(1'b0),.RXDFELFHOLD(1'b0),.RXDFELFOVRDEN(1'b0),.RXDFELPMRESET(1'b0),.RXDFETAP2HOLD(1'b0),.RXDFETAP2OVRDEN(1'b0),.RXDFETAP3HOLD(1'b0),.RXDFETAP3OVRDEN(1'b0),.RXDFETAP4HOLD(1'b0),.RXDFETAP4OVRDEN(1'b0),.RXDFETAP5HOLD(1'b0),.RXDFETAP5OVRDEN(1'b0),.RXDFEUTHOLD(1'b0),.RXDFEUTOVRDEN(1'b0),.RXDFEVPHOLD(1'b0),.RXDFEVPOVRDEN(1'b0),.RXDFEVSEN(1'b0),.RXLPMLFKLOVRDEN(1'b0),.RXMONITOROUT(),.RXMONITORSEL(2'b0),.RXOSHOLD(1'b0),.RXOSOVRDEN(1'b0),.RXRATEDONE(),.RXOUTCLKFABRIC(),.RXOUTCLKPCS(),.RXOUTCLKSEL(3'b010),.RXDATAVALID(),.RXHEADER(),.RXHEADERVALID(),.RXSTARTOFSEQ(),.RXGEARBOXSLIP(1'b0),.RXOOBRESET(1'b0),.RXPCSRESET(1'b0),.RXLPMEN(1'b1),.RXCOMSASDET(),.RXCOMWAKEDET(),.RXCOMINITDET(),.RXELECIDLE(),.RXELECIDLEMODE(2'b11),.RXPOLARITY(1'b0),.RXSLIDE(1'b0),.RXCHBONDI(5'b00000),.RXQPIEN(1'b0),.RXQPISENN(),.RXQPISENP(),.TXPHDLYTSTCLK(1'b0),.TXPOSTCURSOR(5'b0),.TXPOSTCURSORINV(1'b0),.TXPRECURSOR(5'b0),.TXPRECURSORINV(1'b0),.TXQPIBIASEN(1'b0),.TXQPISTRONGPDOWN(1'b0),.TXQPIWEAKPUP(1'b0),.CFGRESET(1'b0),.PCSRSVDOUT(),.GTRESETSEL(1'b0),.RESETOVRD(1'b0),.TXELECIDLE(1'b0),.TXMARGIN(3'b0),.TXRATE(3'b0),.TXSWING(1'b0),.TXPRBSFORCEERR(1'b0),.TXDLYBYPASS(1'b1),.TXDLYEN(1'b0),.TXDLYHOLD(1'b0),.TXDLYOVRDEN(1'b0),.TXDLYSRESET(1'b0),.TXDLYSRESETDONE(),.TXDLYUPDOWN(1'b0),.TXPHALIGN(1'b0),.TXPHALIGNDONE(),.TXPHALIGNEN(1'b0),.TXPHDLYPD(1'b0),.TXPHDLYRESET(1'b0),.TXPHINIT(1'b0),.TXPHINITDONE(),.TXPHOVRDEN(1'b0),.TXBUFSTATUS(),.TXBUFDIFFCTRL(3'b100),.TXDEEMPH(1'b0),.TXDIFFCTRL(4'b1000),.TXDIFFPD(1'b0),.TXINHIBIT(1'b0),.TXMAINCURSOR(7'b0000000),.TXPISOPD(1'b0),.TXOUTCLKFABRIC(),.TXOUTCLKPCS(),.TXOUTCLKSEL(3'b100),.TXRATEDONE(),.TXGEARBOXREADY(),.TXHEADER(3'b0),.TXSEQUENCE(7'b0),.TXSTARTSEQ(1'b0),.TXPCSRESET(1'b0),.TXPMARESET(1'b0),.TXCOMFINISH(),.TXCOMINIT(1'b0),.TXCOMSAS(1'b0),.TXCOMWAKE(1'b0),.TXPDELECIDLEMODE(1'b0),.TXPOLARITY(1'b0),.TXDETECTRX(1'b0),.TX8B10BBYPASS(8'b0),.TXPRBSSEL(3'b0),.TXQPISENN(),.TXQPISENP(),.RXMCOMMAALIGNEN(1'b1),.RXPCOMMAALIGNEN(1'b1),.CPLLPD(1'b0)
,.TXCHARDISPMODE(8'b0)
,.TXCHARDISPVAL({8'b0})
,.CPLLREFCLKSEL
,.RXDISPERR({rxdisperr_float_i,RXDISPERR})
,.RXNOTINTABLE({rxnotintable_float_i,RXNOTINTABLE})
,.RXCHARISCOMMA({rxchariscomma_float_i,RXCHARISCOMMA})
,.RXCHARISK({rxcharisk_float_i,RXCHARISK})
,.TXCHARISK(txcharisk)
,.TXDATA(txdata)
,.RXDATA({rxdata_dummy,RXDATA})
,.GTXTXN,.GTXTXP,.GTXRXP,.GTXRXN,.GTNORTHREFCLK0,.GTNORTHREFCLK1,.GTREFCLK0,.GTREFCLK1,.GTSOUTHREFCLK0,.GTSOUTHREFCLK1,.QPLLCLK,.QPLLREFCLK,.CPLLLOCK,.CPLLRESET,.CPLLFBCLKLOST,.CPLLREFCLKLOST,.CPLLLOCKDETCLK,.RXOUTCLK,.TXOUTCLK,.RXUSRCLK,.RXUSRCLK2,.TXUSRCLK,.TXUSRCLK2,.RXUSERRDY,.RXBYTEISALIGNED,.RXBYTEREALIGN,.RXCOMMADET,.GTRXRESET,.RXPMARESET,.RXRESETDONE,.GTTXRESET,.TXUSERRDY,.TXRESETDONE,.RXVALID
);

wire txclk62_5;
wire txclk62_5_90;
wire txclk125;
wire mmcm_txclkfbout,mmcm_txclkfbin,mmcm_txclk125,mmcm_txclk62_5,mmcm_txclk62_5_90;
MMCME2_BASE #(.BANDWIDTH("OPTIMIZED")
,.CLKIN1_PERIOD(16.0)
,.CLKFBOUT_MULT_F(16)
,.DIVCLK_DIVIDE(1)
,.CLKFBOUT_PHASE(0.0)
,.CLKOUT0_DIVIDE_F(8)
,.CLKOUT0_DUTY_CYCLE(0.5)
,.CLKOUT0_PHASE(0.0)
,.CLKOUT1_DIVIDE(16)
,.CLKOUT1_DUTY_CYCLE(0.5)
,.CLKOUT1_PHASE(0.0)
,.CLKOUT2_DIVIDE(16)
,.CLKOUT2_DUTY_CYCLE(0.5)
,.CLKOUT2_PHASE(90.0)
,.REF_JITTER1(0.0)
,.STARTUP_WAIT("FALSE")
) mmcme2_base_tx(.CLKIN1(mmcm_txoutclk)

,.CLKOUT0(mmcm_txclk125)
,.CLKOUT1(mmcm_txclk62_5)
,.CLKOUT2(mmcm_txclk62_5_90)
,.LOCKED(mmcm_txlocked)
,.CLKFBOUT(mmcm_txclkfbout)
,.CLKFBIN(mmcm_txclkfbin)
,.PWRDWN(1'b0)
,.RST(mmcm_txreset));
BUFG bufgtxoutclk(.I(TXOUTCLK),.O(mmcm_txoutclk));
BUFG mmcmtxclkfb(.I(mmcm_txclkfbout),.O(mmcm_txclkfbin));
BUFG bufgtxclk125(.I(mmcm_txclk125),.O(txclk125));
BUFG bufgtxclk62_5(.I(mmcm_txclk62_5),.O(txclk62_5));
BUFG bufgtxclk62_5_90(.I(mmcm_txclk62_5_90),.O(txclk62_5_90));
assign TXUSRCLK=txclk62_5;
assign TXUSRCLK2=txclk62_5;
assign txusrclk=txclk62_5_90;
assign txusrclk2=txclk125;
wire rxclk62_5;
wire rxclk125;
wire mmcm_rxclkfbout,mmcm_rxclkfbin,mmcm_rxclk125,mmcm_rxclk62_5;
MMCME2_BASE #(.BANDWIDTH("OPTIMIZED"),.CLKIN1_PERIOD(16.0),.CLKFBOUT_MULT_F(16),.DIVCLK_DIVIDE(1),.CLKFBOUT_PHASE(0.0),.CLKOUT0_DIVIDE_F(8),.CLKOUT0_DUTY_CYCLE(0.5),.CLKOUT0_PHASE(0.0),.CLKOUT1_DIVIDE(16),.CLKOUT1_DUTY_CYCLE(0.5),.CLKOUT1_PHASE(0.0),.REF_JITTER1(0.0),.STARTUP_WAIT("FALSE")
) mmcme2_base_rx(.CLKIN1(mmcm_rxoutclk)
,.CLKOUT0(mmcm_rxclk125),.CLKOUT1(mmcm_rxclk62_5),.LOCKED(mmcm_rxlocked),.CLKFBOUT(mmcm_rxclkfbout),.CLKFBIN(mmcm_rxclkfbin),.PWRDWN(1'b0),.RST(mmcm_rxreset));
BUFG bufgrxoutclk(.I(TXOUTCLK),.O(mmcm_rxoutclk));
BUFG mmcmrxclkfb(.I(mmcm_rxclkfbout),.O(mmcm_rxclkfbin));
BUFG bufgrxclk125(.I(mmcm_rxclk125),.O(rxclk125));
BUFG bufgrxclk62_5(.I(mmcm_rxclk62_5),.O(rxclk62_5));
assign RXUSRCLK=rxclk62_5;
assign RXUSRCLK2=rxclk62_5;
assign rxusrclk=rxclk62_5;
assign rxusrclk2=rxclk125;
/*BUFG txoutclk_bufg(.I(TXOUTCLK),.O(TXUSRCLK));
assign TXUSRCLK2=TXUSRCLK;
BUFG rxoutclk_bufg(.I(RXOUTCLK),.O(RXUSRCLK));
assign RXUSRCLK2=RXUSRCLK;
assign txusrclk=TXUSRCLK;
assign rxusrclk=RXUSRCLK;
*/


localparam NSTEP=3;
wire [NSTEP-1:0] done;
wire [NSTEP-1:0] donestrobe;
wire [NSTEP-1:0] error;
wire [NSTEP-1:0] resetout;
assign {CPLLRESET,txrxreset0,txrxreset1}=resetout;
wire [NSTEP-1:0] resetin={reset,donestrobe[NSTEP-1:1]};
wire [NSTEP-1:0] donecriteria={rdyfortxrxreset,txrxresetdone,txrxresetdone};
wire [NSTEP-1:0] readycriteria={readyforreset,donecriteria[NSTEP-1:1],};
wire [NSTEP*16-1:0] readylength={16'd10,16'd10,16'd10};
wire [NSTEP*16-1:0] resetlength={16'd10,16'd10,16'd10};
wire [NSTEP*32-1:0] timeout={NSTEP{32'b0}};
chainreset #(.NSTEP(NSTEP))
chainreset(.clk(CPLLLOCKDETCLK)
,.done,.donecriteria,.donestrobe,.error,.readycriteria,.readylength,.resetin,.resetlength,.resetout,.timeout);
assign resetdone=&done;
assign rdyfortxrxreset=&{readyforreset,CPLLLOCK};
assign txrxresetdone=&{TXRESETDONE,RXRESETDONE,rdyfortxrxreset};
endmodule


