parameter INIT_acqbuf0=""
,parameter INIT_acqbuf1=""
,parameter INIT_command0=""
,parameter INIT_command1=""
,parameter INIT_command2=""
,parameter INIT_command3=""
,parameter INIT_command4=""
,parameter INIT_command5=""
,parameter INIT_command6=""
,parameter INIT_command7=""
,parameter INIT_qdrvfreq0=""
,parameter INIT_qdrvfreq1=""
,parameter INIT_qdrvfreq2=""
,parameter INIT_qdrvfreq3=""
,parameter INIT_qdrvfreq4=""
,parameter INIT_qdrvfreq5=""
,parameter INIT_qdrvfreq6=""
,parameter INIT_qdrvfreq7=""
,parameter INIT_rdrvfreq0=""
,parameter INIT_rdrvfreq1=""
,parameter INIT_rdrvfreq2=""
,parameter INIT_rdrvfreq3=""
,parameter INIT_rdrvfreq4=""
,parameter INIT_rdrvfreq5=""
,parameter INIT_rdrvfreq6=""
,parameter INIT_rdrvfreq7=""
,parameter INIT_dacmon0=""
,parameter INIT_dacmon1=""
,parameter INIT_dacmon2=""
,parameter INIT_dacmon3=""
,parameter INIT_qdrvenv0=""
,parameter INIT_qdrvenv1=""
,parameter INIT_qdrvenv2=""
,parameter INIT_qdrvenv3=""
,parameter INIT_qdrvenv4=""
,parameter INIT_qdrvenv5=""
,parameter INIT_qdrvenv6=""
,parameter INIT_qdrvenv7=""
,parameter INIT_rdloenv0=""
,parameter INIT_rdloenv1=""
,parameter INIT_rdloenv2=""
,parameter INIT_rdloenv3=""
,parameter INIT_rdloenv4=""
,parameter INIT_rdloenv5=""
,parameter INIT_rdloenv6=""
,parameter INIT_rdloenv7=""
,parameter INIT_rdrvenv0=""
,parameter INIT_rdrvenv1=""
,parameter INIT_rdrvenv2=""
,parameter INIT_rdrvenv3=""
,parameter INIT_rdrvenv4=""
,parameter INIT_rdrvenv5=""
,parameter INIT_rdrvenv6=""
,parameter INIT_rdrvenv7=""
,parameter INIT_accbuf0=""
,parameter INIT_accbuf1=""
,parameter INIT_accbuf2=""
,parameter INIT_accbuf3=""
,parameter INIT_accbuf4=""
,parameter INIT_accbuf5=""
,parameter INIT_accbuf6=""
,parameter INIT_accbuf7=""
,parameter INIT_rdlofreq0=""
,parameter INIT_rdlofreq1=""
,parameter INIT_rdlofreq2=""
,parameter INIT_rdlofreq3=""
,parameter INIT_rdlofreq4=""
,parameter INIT_rdlofreq5=""
,parameter INIT_rdlofreq6=""
,parameter INIT_rdlofreq7=""
,parameter INIT_sdbuf0=""
,parameter INIT_sdbuf1=""
,parameter INIT_sdbuf2=""
,parameter INIT_sdbuf3=""
,parameter INIT_sdbuf4=""
,parameter INIT_sdbuf5=""
,parameter INIT_sdbuf6=""
,parameter INIT_sdbuf7=""
,parameter INIT_sdpara0=""
,parameter INIT_sdpara1=""
,parameter INIT_sdpara2=""
,parameter INIT_sdpara3=""
,parameter INIT_sdpara4=""
,parameter INIT_sdpara5=""
,parameter INIT_sdpara6=""
,parameter INIT_sdpara7=""