.acqbuf0_R(acqbuf0_R)
,.acqbuf1_R(acqbuf1_R)
,.command0_W(command0_W)
,.command1_W(command1_W)
,.command2_W(command2_W)
,.command3_W(command3_W)
,.command4_W(command4_W)
,.command5_W(command5_W)
,.command6_W(command6_W)
,.command7_W(command7_W)
,.qdrvfreq0_W(qdrvfreq0_W)
,.qdrvfreq1_W(qdrvfreq1_W)
,.qdrvfreq2_W(qdrvfreq2_W)
,.qdrvfreq3_W(qdrvfreq3_W)
,.qdrvfreq4_W(qdrvfreq4_W)
,.qdrvfreq5_W(qdrvfreq5_W)
,.qdrvfreq6_W(qdrvfreq6_W)
,.qdrvfreq7_W(qdrvfreq7_W)
,.rdrvfreq0_W(rdrvfreq0_W)
,.rdrvfreq1_W(rdrvfreq1_W)
,.rdrvfreq2_W(rdrvfreq2_W)
,.rdrvfreq3_W(rdrvfreq3_W)
,.rdrvfreq4_W(rdrvfreq4_W)
,.rdrvfreq5_W(rdrvfreq5_W)
,.rdrvfreq6_W(rdrvfreq6_W)
,.rdrvfreq7_W(rdrvfreq7_W)
,.dacmon0_R(dacmon0_R)
,.dacmon1_R(dacmon1_R)
,.dacmon2_R(dacmon2_R)
,.dacmon3_R(dacmon3_R)
,.qdrvenv0_W(qdrvenv0_W)
,.qdrvenv1_W(qdrvenv1_W)
,.qdrvenv2_W(qdrvenv2_W)
,.qdrvenv3_W(qdrvenv3_W)
,.qdrvenv4_W(qdrvenv4_W)
,.qdrvenv5_W(qdrvenv5_W)
,.qdrvenv6_W(qdrvenv6_W)
,.qdrvenv7_W(qdrvenv7_W)
,.rdloenv0_W(rdloenv0_W)
,.rdloenv1_W(rdloenv1_W)
,.rdloenv2_W(rdloenv2_W)
,.rdloenv3_W(rdloenv3_W)
,.rdloenv4_W(rdloenv4_W)
,.rdloenv5_W(rdloenv5_W)
,.rdloenv6_W(rdloenv6_W)
,.rdloenv7_W(rdloenv7_W)
,.rdrvenv0_W(rdrvenv0_W)
,.rdrvenv1_W(rdrvenv1_W)
,.rdrvenv2_W(rdrvenv2_W)
,.rdrvenv3_W(rdrvenv3_W)
,.rdrvenv4_W(rdrvenv4_W)
,.rdrvenv5_W(rdrvenv5_W)
,.rdrvenv6_W(rdrvenv6_W)
,.rdrvenv7_W(rdrvenv7_W)
,.accbuf0_R(accbuf0_R)
,.accbuf1_R(accbuf1_R)
,.accbuf2_R(accbuf2_R)
,.accbuf3_R(accbuf3_R)
,.accbuf4_R(accbuf4_R)
,.accbuf5_R(accbuf5_R)
,.accbuf6_R(accbuf6_R)
,.accbuf7_R(accbuf7_R)
,.rdlofreq0_W(rdlofreq0_W)
,.rdlofreq1_W(rdlofreq1_W)
,.rdlofreq2_W(rdlofreq2_W)
,.rdlofreq3_W(rdlofreq3_W)
,.rdlofreq4_W(rdlofreq4_W)
,.rdlofreq5_W(rdlofreq5_W)
,.rdlofreq6_W(rdlofreq6_W)
,.rdlofreq7_W(rdlofreq7_W)
,.sdbuf0_R(sdbuf0_R)
,.sdbuf1_R(sdbuf1_R)
,.sdbuf2_R(sdbuf2_R)
,.sdbuf3_R(sdbuf3_R)
,.sdbuf4_R(sdbuf4_R)
,.sdbuf5_R(sdbuf5_R)
,.sdbuf6_R(sdbuf6_R)
,.sdbuf7_R(sdbuf7_R)