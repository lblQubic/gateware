wire DAC00_M_AXIS_ACLK;
    wire DAC00_M_AXIS_ARESETN;
    wire  DAC00_M_AXIS_TREADY;
    wire  DAC00_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC00_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC00_M_AXIS_TSTRB;
    wire  DAC00_M_AXIS_TLAST;
    
wire DAC01_M_AXIS_ACLK;
    wire DAC01_M_AXIS_ARESETN;
    wire  DAC01_M_AXIS_TREADY;
    wire  DAC01_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC01_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC01_M_AXIS_TSTRB;
    wire  DAC01_M_AXIS_TLAST;
    
wire DAC02_M_AXIS_ACLK;
    wire DAC02_M_AXIS_ARESETN;
    wire  DAC02_M_AXIS_TREADY;
    wire  DAC02_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC02_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC02_M_AXIS_TSTRB;
    wire  DAC02_M_AXIS_TLAST;
    
wire DAC03_M_AXIS_ACLK;
    wire DAC03_M_AXIS_ARESETN;
    wire  DAC03_M_AXIS_TREADY;
    wire  DAC03_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC03_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC03_M_AXIS_TSTRB;
    wire  DAC03_M_AXIS_TLAST;
    
wire DAC10_M_AXIS_ACLK;
    wire DAC10_M_AXIS_ARESETN;
    wire  DAC10_M_AXIS_TREADY;
    wire  DAC10_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC10_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC10_M_AXIS_TSTRB;
    wire  DAC10_M_AXIS_TLAST;
    
wire DAC11_M_AXIS_ACLK;
    wire DAC11_M_AXIS_ARESETN;
    wire  DAC11_M_AXIS_TREADY;
    wire  DAC11_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC11_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC11_M_AXIS_TSTRB;
    wire  DAC11_M_AXIS_TLAST;
    
wire DAC12_M_AXIS_ACLK;
    wire DAC12_M_AXIS_ARESETN;
    wire  DAC12_M_AXIS_TREADY;
    wire  DAC12_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC12_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC12_M_AXIS_TSTRB;
    wire  DAC12_M_AXIS_TLAST;
    
wire DAC13_M_AXIS_ACLK;
    wire DAC13_M_AXIS_ARESETN;
    wire  DAC13_M_AXIS_TREADY;
    wire  DAC13_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC13_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC13_M_AXIS_TSTRB;
    wire  DAC13_M_AXIS_TLAST;
    
wire DAC20_M_AXIS_ACLK;
    wire DAC20_M_AXIS_ARESETN;
    wire  DAC20_M_AXIS_TREADY;
    wire  DAC20_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC20_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC20_M_AXIS_TSTRB;
    wire  DAC20_M_AXIS_TLAST;
    
wire DAC21_M_AXIS_ACLK;
    wire DAC21_M_AXIS_ARESETN;
    wire  DAC21_M_AXIS_TREADY;
    wire  DAC21_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC21_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC21_M_AXIS_TSTRB;
    wire  DAC21_M_AXIS_TLAST;
    
wire DAC22_M_AXIS_ACLK;
    wire DAC22_M_AXIS_ARESETN;
    wire  DAC22_M_AXIS_TREADY;
    wire  DAC22_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC22_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC22_M_AXIS_TSTRB;
    wire  DAC22_M_AXIS_TLAST;
    
wire DAC23_M_AXIS_ACLK;
    wire DAC23_M_AXIS_ARESETN;
    wire  DAC23_M_AXIS_TREADY;
    wire  DAC23_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC23_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC23_M_AXIS_TSTRB;
    wire  DAC23_M_AXIS_TLAST;
    
wire DAC30_M_AXIS_ACLK;
    wire DAC30_M_AXIS_ARESETN;
    wire  DAC30_M_AXIS_TREADY;
    wire  DAC30_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC30_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC30_M_AXIS_TSTRB;
    wire  DAC30_M_AXIS_TLAST;
    
wire DAC31_M_AXIS_ACLK;
    wire DAC31_M_AXIS_ARESETN;
    wire  DAC31_M_AXIS_TREADY;
    wire  DAC31_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC31_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC31_M_AXIS_TSTRB;
    wire  DAC31_M_AXIS_TLAST;
    
wire DAC32_M_AXIS_ACLK;
    wire DAC32_M_AXIS_ARESETN;
    wire  DAC32_M_AXIS_TREADY;
    wire  DAC32_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC32_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC32_M_AXIS_TSTRB;
    wire  DAC32_M_AXIS_TLAST;
    
wire DAC33_M_AXIS_ACLK;
    wire DAC33_M_AXIS_ARESETN;
    wire  DAC33_M_AXIS_TREADY;
    wire  DAC33_M_AXIS_TVALID;
    wire  [DAC_AXIS_DATAWIDTH-1 : 0] DAC33_M_AXIS_TDATA;
    wire  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC33_M_AXIS_TSTRB;
    wire  DAC33_M_AXIS_TLAST;
    
wire  ADC00_S_AXIS_ACLK;
    wire  ADC00_S_AXIS_ARESETN;
    wire  ADC00_S_AXIS_TREADY;
    wire  ADC00_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC00_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC00_S_AXIS_TSTRB;
    wire  ADC00_S_AXIS_TLAST;
    
wire  ADC01_S_AXIS_ACLK;
    wire  ADC01_S_AXIS_ARESETN;
    wire  ADC01_S_AXIS_TREADY;
    wire  ADC01_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC01_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC01_S_AXIS_TSTRB;
    wire  ADC01_S_AXIS_TLAST;
    
wire  ADC02_S_AXIS_ACLK;
    wire  ADC02_S_AXIS_ARESETN;
    wire  ADC02_S_AXIS_TREADY;
    wire  ADC02_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC02_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC02_S_AXIS_TSTRB;
    wire  ADC02_S_AXIS_TLAST;
    
wire  ADC03_S_AXIS_ACLK;
    wire  ADC03_S_AXIS_ARESETN;
    wire  ADC03_S_AXIS_TREADY;
    wire  ADC03_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC03_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC03_S_AXIS_TSTRB;
    wire  ADC03_S_AXIS_TLAST;
    
wire  ADC10_S_AXIS_ACLK;
    wire  ADC10_S_AXIS_ARESETN;
    wire  ADC10_S_AXIS_TREADY;
    wire  ADC10_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC10_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC10_S_AXIS_TSTRB;
    wire  ADC10_S_AXIS_TLAST;
    
wire  ADC11_S_AXIS_ACLK;
    wire  ADC11_S_AXIS_ARESETN;
    wire  ADC11_S_AXIS_TREADY;
    wire  ADC11_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC11_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC11_S_AXIS_TSTRB;
    wire  ADC11_S_AXIS_TLAST;
    
wire  ADC12_S_AXIS_ACLK;
    wire  ADC12_S_AXIS_ARESETN;
    wire  ADC12_S_AXIS_TREADY;
    wire  ADC12_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC12_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC12_S_AXIS_TSTRB;
    wire  ADC12_S_AXIS_TLAST;
    
wire  ADC13_S_AXIS_ACLK;
    wire  ADC13_S_AXIS_ARESETN;
    wire  ADC13_S_AXIS_TREADY;
    wire  ADC13_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC13_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC13_S_AXIS_TSTRB;
    wire  ADC13_S_AXIS_TLAST;
    
wire  ADC20_S_AXIS_ACLK;
    wire  ADC20_S_AXIS_ARESETN;
    wire  ADC20_S_AXIS_TREADY;
    wire  ADC20_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC20_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC20_S_AXIS_TSTRB;
    wire  ADC20_S_AXIS_TLAST;
    
wire  ADC21_S_AXIS_ACLK;
    wire  ADC21_S_AXIS_ARESETN;
    wire  ADC21_S_AXIS_TREADY;
    wire  ADC21_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC21_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC21_S_AXIS_TSTRB;
    wire  ADC21_S_AXIS_TLAST;
    
wire  ADC22_S_AXIS_ACLK;
    wire  ADC22_S_AXIS_ARESETN;
    wire  ADC22_S_AXIS_TREADY;
    wire  ADC22_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC22_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC22_S_AXIS_TSTRB;
    wire  ADC22_S_AXIS_TLAST;
    
wire  ADC23_S_AXIS_ACLK;
    wire  ADC23_S_AXIS_ARESETN;
    wire  ADC23_S_AXIS_TREADY;
    wire  ADC23_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC23_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC23_S_AXIS_TSTRB;
    wire  ADC23_S_AXIS_TLAST;
    
wire  ADC30_S_AXIS_ACLK;
    wire  ADC30_S_AXIS_ARESETN;
    wire  ADC30_S_AXIS_TREADY;
    wire  ADC30_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC30_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC30_S_AXIS_TSTRB;
    wire  ADC30_S_AXIS_TLAST;
    
wire  ADC31_S_AXIS_ACLK;
    wire  ADC31_S_AXIS_ARESETN;
    wire  ADC31_S_AXIS_TREADY;
    wire  ADC31_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC31_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC31_S_AXIS_TSTRB;
    wire  ADC31_S_AXIS_TLAST;
    
wire  ADC32_S_AXIS_ACLK;
    wire  ADC32_S_AXIS_ARESETN;
    wire  ADC32_S_AXIS_TREADY;
    wire  ADC32_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC32_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC32_S_AXIS_TSTRB;
    wire  ADC32_S_AXIS_TLAST;
    
wire  ADC33_S_AXIS_ACLK;
    wire  ADC33_S_AXIS_ARESETN;
    wire  ADC33_S_AXIS_TREADY;
    wire  ADC33_S_AXIS_TVALID;
    wire  [ADC_AXIS_DATAWIDTH-1 : 0] ADC33_S_AXIS_TDATA;
    wire  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC33_S_AXIS_TSTRB;
    wire  ADC33_S_AXIS_TLAST;
    