module boardcfg #(
`include "plps_para.vh"	
,`include "bram_para.vh"
,`include "braminit_para.vh"
)(hwif.cfg hw
,ifcfgregs.regs cfgregs
,ifdspregs.regs dspregs
,`include "bramif_port.vh"
,`include "rfdcif_port.vh"
,ifdsp.cfg dspif
,output cfgclk
,output dspclk
,input pl_clk0
,input clk_dac0
,input clk_dac1
,input clk_dac2
,input clk_dac3
,input clk_adc0
,input clk_adc1
,input clk_adc2
,input clk_adc3
,input clkadc3_300
,input clkadc3_600
,input aresetn
,output cfgreset
,output dspreset
,output psreset
,output adc3reset
);
wire reset=(~aresetn)|hw.gpio_sw_c;
areset #(.WIDTH(1),.SRWIDTH(4))
cfgareset(.clk(cfgclk),.areset(reset),.sreset(cfgreset),.sreset_val());
areset #(.WIDTH(1),.SRWIDTH(4))
dspareset(.clk(dspclk),.areset(reset),.sreset(dspreset),.sreset_val());
areset #(.WIDTH(1),.SRWIDTH(4))
psareset(.clk(pl_clk0),.areset(reset),.sreset(psreset),.sreset_val());
areset #(.WIDTH(1),.SRWIDTH(4))
adc3areset(.clk(clkadc3_600),.areset(reset),.sreset(adc3reset),.sreset_val());

gitrevision gitrevision(cfgregs.gitrevision);


reg [31:0] cnt100=0;
always @(posedge hw.clk100) begin
	cnt100<=cnt100+1;
end
reg [31:0] cnt125=0;
always @(posedge hw.clk125) begin
	cnt125<=cnt125+1;
end
assign cfgclk=hw.clk100;
assign dspclk=hw.clk104_pl_clk;// clk_dac2;
//assign dspclk=clk_dac2;
assign hw.ledrgb[0][1]=cnt100[27];
assign hw.ledrgb[1][1]=cnt100[26];
assign hw.ledrgb[2][1]=cnt100[25];
assign hw.ledrgb[3][1]=cnt100[24];

assign hw.ledrgb[4][1]=cnt125[27];
assign hw.ledrgb[5][1]=cnt125[26];
assign hw.ledrgb[6][1]=cnt125[25];
assign hw.ledrgb[7][1]=cnt125[24];

//assign regs.test1=regs.r0+regs.r1+regs.r2+regs.r3;
assign hw.ledrgb[0][0]=cfgregs.test1[0];
assign hw.ledrgb[1][0]=cfgregs.test1[1];
assign hw.ledrgb[2][0]=cfgregs.test1[2];
assign hw.ledrgb[3][0]=cfgregs.test1[3];
assign hw.ledrgb[4][0]=cfgregs.test1[4];
assign hw.ledrgb[5][0]=cfgregs.test1[5];
assign hw.ledrgb[6][0]=cfgregs.test1[6];
assign hw.ledrgb[7][0]=cfgregs.test1[7];
/*assign hw.pmod0[6]=cnt100[1];
assign hw.pmod0[5]=cnt125[1];
assign hw.pmod0[4]=hw.usersi570c0;
assign hw.pmod0[3]=hw.usersi570c1;
assign hw.pmod0[2]=hw.clk104_pl_sysref;
assign hw.pmod0[1]=hw.clk104_pl_clk;
*/
assign hw.ledrgb[0][2]=cfgregs.test[0];
assign hw.ledrgb[1][2]=cfgregs.test[1];
assign hw.ledrgb[2][2]=cfgregs.test[2];
assign hw.ledrgb[3][2]=cfgregs.test[3];
assign hw.ledrgb[4][2]=cfgregs.test[4];
assign hw.ledrgb[5][2]=cfgregs.test[5];
assign hw.ledrgb[6][2]=cfgregs.test[6];
assign hw.ledrgb[7][2]=cfgregs.test[7];

enum {CLK100
,CLK125
,USERSI570C0
,USERSI570C1
,CLK104PLSYSREF
,CLK104PLCLK
,CLKDAC0
,CLKDAC1
,CLKDAC2
,CLKDAC3
,CLKADC0
,CLKADC1
,CLKADC2
,CLKADC3
,CLKADC3_300
,CLKADC3_600
//,MGTREFCLK1_X0Y1
,NFCNT
} fcnt;

wire [32*NFCNT-1:0] freq_cnt;
assign freq_cnt={cfgregs.fclk100
,cfgregs.fclk125
,cfgregs.fusersi570c0
,cfgregs.fusersi570c1
,cfgregs.fclk104plsysref
,cfgregs.fclk104plclk
,cfgregs.fclk_dac0
,cfgregs.fclk_dac1
,cfgregs.fclk_dac2
,cfgregs.fclk_dac3
,cfgregs.fclk_adc0
,cfgregs.fclk_adc1
,cfgregs.fclk_adc2
,cfgregs.fclk_adc3
,cfgregs.fclkadc3_300
,cfgregs.fclkadc3_600
};

wire [NFCNT-1:0] freqcnt_clks= {
	hw.clk100
	,hw.clk125
	,hw.usersi570c0
	,hw.usersi570c1
	,hw.clk104_pl_sysref
	,hw.clk104_pl_clk
	,clk_dac0
	,clk_dac1
	,clk_dac2
	,clk_dac3
	,clk_adc0
	,clk_adc1
	,clk_adc2
	,clk_adc3
	,clkadc3_300
	,clkadc3_600
};

genvar jx;
generate for (jx=0; jx<NFCNT; jx=jx+1)	begin: gen_fcnt
	freq_count3 #(.REFCNTWIDTH(24))
	freq_count3(.clk(hw.clk100),.fin(freqcnt_clks[jx]),.frequency(freq_cnt[jx*32+31:jx*32]));
//		{regs.fclk100,regs.fclk125,regs.fusersi570c0,regs.fusersi570c1,regs.fclk104plsysref,regs.fclk104plclk,regs.fclk_dac2,regs.fclk_dac3,regs.fclk_adc2,regs.fclkadc2_300,regs.fclkadc2_600}
end
endgenerate

`include "bram_read.vh"
`include "bram_write.vh"

//wire adc00datavalid;
//axi4stream_slave_handshake_data #(.DATA_WIDTH (ADC_AXIS_DATAWIDTH))adc00hsda(.axis(adc00axis),.ready(1'b1),.datavalid(adc00datavalid),.data(dspif.adc[0]));
//wire adc20datavalid;
//axi4stream_slave_handshake_data #(.DATA_WIDTH (ADC_AXIS_DATAWIDTH))adc20hsda(.axis(adc20axis),.ready(1'b1),.datavalid(adc20datavalid),.data(dspif.adc[1]));
wire adc30datavalid;
axi4stream_slave_handshake_data #(.DATA_WIDTH (ADC_AXIS_DATAWIDTH))adc30hsda(.axis(adc30axis),.ready(1'b1),.datavalid(adc30datavalid),.data(dspif.adc[1]));
wire adc32datavalid;
axi4stream_slave_handshake_data #(.DATA_WIDTH (ADC_AXIS_DATAWIDTH))adc32hsda(.axis(adc32axis),.ready(1'b1),.datavalid(adc32datavalid),.data(dspif.adc[0]));

axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac00hsda(.axis(dac00axis),.datavalid(1'b1),.data(dspif.dac[8])); // 228 0
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac01hsda(.axis(dac01axis),.datavalid(1'b1),.data(dspif.dac[3])); // 228 1
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac02hsda(.axis(dac02axis),.datavalid(1'b1),.data(dspif.dac[2])); // 228 2
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac03hsda(.axis(dac03axis),.datavalid(1'b1),.data(dspif.dac[4])); // 228 3
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac10hsda(.axis(dac10axis),.datavalid(1'b1),.data(dspif.dac[1])); // 229 0
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac11hsda(.axis(dac11axis),.datavalid(1'b1),.data(dspif.dac[5])); // 229 1
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac12hsda(.axis(dac12axis),.datavalid(1'b1),.data(dspif.dac[0])); // 229 2
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac13hsda(.axis(dac13axis),.datavalid(1'b1),.data(dspif.dac[6])); // 229 3
axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac20hsda(.axis(dac20axis),.datavalid(1'b1),.data(dspif.dac[7])); // 230 0
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac21hsda(.axis(dac21axis),.datavalid(1'b1),.data(dspif.dac[9]));
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac22hsda(.axis(dac22axis),.datavalid(1'b1),.data(dspif.dac[10]));
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac23hsda(.axis(dac23axis),.datavalid(1'b1),.data(dspif.dac[11]));
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac30hsda(.axis(dac30axis),.datavalid(1'b1),.data(dspif.dac[12]));
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac31hsda(.axis(dac31axis),.datavalid(1'b1),.data(dspif.dac[13]));
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac32hsda(.axis(dac32axis),.datavalid(1'b1),.data(dspif.dac[14]));
//axi4stream_master_handshake_data #(.DATA_WIDTH (DAC_AXIS_DATAWIDTH))dac33hsda(.axis(dac33axis),.datavalid(1'b1),.data(dspif.dac[15]));
//assign dspif.clk=dspclk;
reg dspreset_r=0;
always @(posedge dspclk) begin
	dspreset_r<=dspreset|dspregs.wstb_dspreset;
end
assign dspif.reset=dspreset_r;

assign dspif.stb_start=dspregs.wstb_start;
assign dspif.start=ready_dspclk;
assign dspif.nshot=dspregs.nshot;
assign dspif.resetacc=dspregs.resetacc;
assign dspif.stb_reset_bram_read=dspregs.wstb_reset_bram_read;
assign dspregs.lastshotdone=dspif.lastshotdone;
assign dspregs.shotcnt=dspif.shotcnt;
assign dspregs.addr_accbuf_mon0=dspif.addr_accbuf_mon0;
assign dspregs.addr_accbuf_mon1=dspif.addr_accbuf_mon1;
assign dspregs.addr_accbuf_mon2=dspif.addr_accbuf_mon2;
assign dspregs.addr_accbuf_mon3=dspif.addr_accbuf_mon3;

assign dspif.acqbufreset=dspregs.acqbufreset;
assign dspif.dacmonreset=dspregs.dacmonreset;
assign dspif.delayaftertrig=dspregs.delayaftertrig;
assign dspif.decimator=dspregs.decimator;
assign dspif.acqchansel[0]=dspregs.acqchansel0;
assign dspif.acqchansel[1]=dspregs.acqchansel1;
assign dspif.dacmonchansel[0]=dspregs.dacmonchansel0;
assign dspif.dacmonchansel[1]=dspregs.dacmonchansel1;
assign dspif.dacmonchansel[2]=dspregs.dacmonchansel2;
assign dspif.dacmonchansel[3]=dspregs.dacmonchansel3;

assign dspif.mixbb1sel=dspregs.mixbb1sel;
assign dspif.mixbb2sel=dspregs.mixbb2sel;
assign dspif.shift=dspregs.shift;


reg current_sample=1'b0;
reg last_sample=1'b0;
reg [2:0] sysref_cnt=0;
reg ready_sysref=1'b0;
always @(posedge dspclk) begin
    current_sample <= hw.clk104_pl_sysref;
    last_sample <= current_sample;
    if (dspregs.start) begin
        sysref_cnt <= sysref_cnt + (~last_sample & current_sample);
    end
    if (sysref_cnt[2]) ready_sysref<=1'b1;
end

assign dspif.test_amp=dspregs.test_amp;
assign dspif.test_freq=dspregs.test_freq;

reg [63:0] dspclkcnt_orig=0;
wire [63:0] corr64={dspregs.copper_corr64_h,dspregs.copper_corr64_l};
reg [63:0] dspclkcnt_corr=0;
always @(posedge dspclk) begin
	if (ready_sysref) dspclkcnt_orig <= dspclkcnt_orig + 1;
	dspclkcnt_corr <= dspclkcnt_orig + corr64;
end

wire dspclkcnt_sw=dspregs.copper_clkcnt_sw;
wire [63:0] dspclkcnt;
assign dspclkcnt = dspclkcnt_sw ? dspclkcnt_corr : dspclkcnt_orig;

wire [63:0] dspclkcnt_trig={dspregs.copper_clkcnt_trig_h,dspregs.copper_clkcnt_trig_l};
reg ready_dspclk=1'b0;
always @(posedge dspclk) begin
	ready_dspclk <= dspclkcnt>=dspclkcnt_trig;
end

// Multi-FPGA synchronization //
wire [63:0] copper_tx_clkcnt;
wire [63:0] copper_rx_clkcnt;
reg [63:0] copper_tx_clkcnt_r=0;
reg [63:0] copper_rx_clkcnt_r=0;
wire copper_tx_data;
wire copper_rx_data;
wire copper_tx_en=dspregs.copper_tx_en;
wire copper_tx_rst=dspregs.copper_tx_rst;

//IOBUF synciobuf (.IO(hw.pmod1[0]),.I(copper_tx_data),.O(copper_rx_data),.T(~copper_tx_en));
IOBUF synciobuf (.IO(hw.dacio[0]),.I(copper_tx_data),.O(copper_rx_data),.T(~copper_tx_en));

//assign hw.pmod1[0]= ~copper_tx_en ? copper_tx_data : 1'bz;
//assign copper_rx_data = hw.pmod1[0];

sync sync_copper(.clk(dspclk)
,.tx_data(copper_tx_data)
,.tx_rst(copper_tx_rst)
,.rx_data(copper_rx_data)
,.clkcnt(dspclkcnt)
,.tx_clkcnt(copper_tx_clkcnt)
,.rx_clkcnt(copper_rx_clkcnt)
);
always @(posedge dspclk) begin
	copper_tx_clkcnt_r<=copper_tx_clkcnt;
	copper_rx_clkcnt_r<=copper_rx_clkcnt;
end
assign	{dspregs.copper_tx_clkcnt_h,dspregs.copper_tx_clkcnt_l}=copper_tx_clkcnt_r;
assign	{dspregs.copper_rx_clkcnt_h,dspregs.copper_rx_clkcnt_l}=copper_rx_clkcnt_r;

// loop back //
wire [63:0] copper_tx_clkcnt_slv;
wire [63:0] copper_rx_clkcnt_slv;
reg [63:0] copper_tx_clkcnt_slv_r=0;
reg [63:0] copper_rx_clkcnt_slv_r=0;
wire copper_tx_data_slv;
wire copper_rx_data_slv;
wire copper_tx_en_slv=dspregs.copper_tx_en_slv;
wire copper_tx_rst_slv=dspregs.copper_tx_rst_slv;

//IOBUF synciobuf_slv (.IO(hw.pmod1[1]),.I(copper_tx_data_slv),.O(copper_rx_data_slv),.T(~copper_tx_en_slv));
IOBUF synciobuf_slv (.IO(hw.dacio[1]),.I(copper_tx_data_slv),.O(copper_rx_data_slv),.T(~copper_tx_en_slv));
//assign hw.pmod1[1]= ~copper_tx_en_slv ? copper_tx_data_slv : 1'bz;
//assign copper_rx_data_slv = hw.pmod1[1];
sync sync_copper_slv(.clk(dspclk)
,.tx_data(copper_tx_data_slv)
,.tx_rst(copper_tx_rst_slv)
,.rx_data(copper_rx_data_slv)
,.clkcnt(dspclkcnt)
,.tx_clkcnt(copper_tx_clkcnt_slv)
,.rx_clkcnt(copper_rx_clkcnt_slv)
);
always @(posedge dspclk) begin
	copper_tx_clkcnt_slv_r<=copper_tx_clkcnt_slv;
	copper_rx_clkcnt_slv_r<=copper_rx_clkcnt_slv;
end
assign	{dspregs.copper_tx_clkcnt_h_slv,dspregs.copper_tx_clkcnt_l_slv}=copper_tx_clkcnt_slv_r;
assign	{dspregs.copper_rx_clkcnt_h_slv,dspregs.copper_rx_clkcnt_l_slv}=copper_rx_clkcnt_slv_r;

//assign hw.pmod1[7:2]=dspclkcnt[25:20];
assign hw.dacio[15:2]=dspclkcnt[25:12];


reg [31:0] coef[0:7][0:7];

wire [31:0] coefused00=dspif.coefused[0][0];
wire [31:0] coefused01=dspif.coefused[0][1];
wire [31:0] coefused02=dspif.coefused[0][2];
wire [31:0] coefused03=dspif.coefused[0][3];
wire [31:0] coefused04=dspif.coefused[0][4];
wire [31:0] coefused05=dspif.coefused[0][5];
wire [31:0] coefused06=dspif.coefused[0][6];
wire [31:0] coefused07=dspif.coefused[0][7];
wire [31:0] coefused10=dspif.coefused[1][0];
wire [31:0] coefused11=dspif.coefused[1][1];
wire [31:0] coefused12=dspif.coefused[1][2];
wire [31:0] coefused13=dspif.coefused[1][3];
wire [31:0] coefused14=dspif.coefused[1][4];
wire [31:0] coefused15=dspif.coefused[1][5];
wire [31:0] coefused16=dspif.coefused[1][6];
wire [31:0] coefused17=dspif.coefused[1][7];
generate
for (genvar i=0;i<8;i=i+1) begin
    for (genvar j=0;j<8;j=j+1) begin
        always @(posedge dspclk) begin
            if (dspregs.wstb_coef) begin
                if (dspregs.waddr_coef==i*8+j) begin
                    dspif.coef[i][j]<=dspregs.wdata_coef;
                end
            end
            if (dspregs.rstb_coefused) begin
                if (dspregs.raddr_coefused==i*8+j) begin
                    dspregs.rdata_coefused<=dspif.coefused[i][j];
                end
            end
        end
    end
end
endgenerate

assign dspregs.procdone=dspif.procdone;
assign dspregs.cnt00=dac00axis.cnt;
assign dspregs.cnt01=dac01axis.cnt;
assign dspregs.cnt02=dac02axis.cnt;
assign dspregs.cnt03=dac03axis.cnt;
assign dspregs.cnt10=dac10axis.cnt;
assign dspregs.cnt11=dac11axis.cnt;
assign dspregs.cnt12=dac12axis.cnt;
assign dspregs.cnt13=dac13axis.cnt;
assign dspregs.cnt20=dac20axis.cnt;

//`include "ilaauto.vh"



wire gtyrxp, gtyrxn;
assign gtyrxp= hw.sfp0_rx_p;
assign gtyrxn= hw.sfp0_rx_n;
wire gtytxp, gtytxn;
assign hw.sfp0_tx_p = gtytxp;
assign hw.sfp0_tx_n = gtytxn;
wire gtwiz_reset_clk_freerun_in;
assign gtwiz_reset_clk_freerun_in = hw.clk125;
wire gtwiz_reset;
assign gtwiz_reset = dspregs.gtwiz_reset;
//assign dspregs.gtwiz_rxdata = gtwiz_userdata_rx;
//assign dspregs.gtwiz_rxctrl0 = rxctrl0;
//assign dspregs.gtwiz_rxctrl1 = rxctrl1;
//assign dspregs.gtwiz_rxctrl2 = rxctrl2;
//assign dspregs.gtwiz_rxctrl3 = rxctrl3;
//assign dspregs.gtwiz_userclk_rx_active = gtwiz_userclk_rx_active;
//assign dspregs.gtwiz_userclk_rx_usrclk2 = gtwiz_userclk_rx_usrclk2;

data_xdomain #(.DWIDTH(32)) usrrx_x_dsp_rxdata (.clkin(gtwiz_userclk_rx_usrclk2),.clkout(dspclk),.gatein(1'b1),.datain(gtwiz_userdata_rx),.gateout(),.dataout(dspregs.gtwiz_rxdata));
data_xdomain #(.DWIDTH(1)) usrrx_x_dsp_rxactive (.clkin(gtwiz_userclk_rx_usrclk2),.clkout(dspclk),.gatein(1'b1),.datain(gtwiz_userclk_rx_active),.gateout(),.dataout(dspregs.gtwiz_userclk_rx_active));

wire gtwiz_reset_all_init;
wire gtwiz_reset_all_buf;
IBUF ibuf_gtwiz_reset_all (.I(gtwiz_reset),.O(gtwiz_reset_all_buf));
wire gtwiz_reset_all;
assign gtwiz_reset_all = gtwiz_reset_all_buf || gtwiz_reset_all_init;

wire gtwiz_reset_clk_freerun_buf;
BUFG bufg_gtwiz_clk_freerun (.I(gtwiz_reset_clk_freerun_in),.O(gtwiz_reset_clk_freerun_buf));

assign gtrefclk00 = hw.mgtrefclk1_128;
assign hw.mgtrefclk0_128= rxrecclkout;

wire gtwiz_userclk_tx_reset;
wire gtwiz_userclk_rx_reset;
assign gtwiz_userclk_tx_reset = ~(&txpmaresetdone);
assign gtwiz_userclk_rx_reset = ~(&rxpmaresetdone);


wire [31:0] gtwiz_txdata;
reg [31:0] dspregs_gtwiz_txdata=0;
always @(posedge dspclk) begin
	dspregs_gtwiz_txdata <= dspregs.gtwiz_txdata;
end
data_xdomain #(.DWIDTH(32)) dsp_x_usrtx_txdata (.clkin(dspclk),.clkout(gtwiz_userclk_tx_usrclk2),.gatein(1'b1),.datain(dspregs_gtwiz_txdata),.gateout(),.dataout(gtwiz_txdata));
//data_xdomain #(.DWIDTH(32)) dsp_x_usrtx_txdata (.clkin(dspclk),.clkout(gtwiz_userclk_tx_usrclk2),.gatein(1'b1),.datain(dspregs.gtwiz_txdata),.gateout(),.dataout(gtwiz_txdata));

gty_sfp_stimulus_8b10b stimulus_inst (
  .gtwiz_reset_all_in          (gtwiz_reset_all || ~gtwiz_reset_rx_done),
  .gtwiz_userclk_tx_usrclk2_in (gtwiz_userclk_tx_usrclk2),
  .gtwiz_userclk_tx_active_in  (gtwiz_userclk_tx_active),
  .txdata_in                   (gtwiz_txdata),
  .txctrl0_out                 (txctrl0),
  .txctrl1_out                 (txctrl1),
  .txctrl2_out                 (txctrl2),
  .txdata_out                  (gtwiz_userdata_tx)
);


wire gtwiz_init_done;
wire [3:0] gtwiz_init_retry_ctr;

wire gtwiz_reset_rx_datapath_init;
assign gtwiz_reset_rx_datapath = gtwiz_reset_rx_datapath_init;

reg gtwiz_sm_link = 1'b1;
gty_sfp_init init_inst (
  .clk_freerun_in  (gtwiz_reset_clk_freerun_buf),
  .reset_all_in    (gtwiz_reset_all),
  .tx_init_done_in (gtwiz_reset_tx_done),
  .rx_init_done_in (gtwiz_reset_rx_done),
  .rx_data_good_in (gtwiz_sm_link),
  .reset_all_out   (gtwiz_reset_all_init),
  .reset_rx_out    (gtwiz_reset_rx_datapath_init),
  .init_done_out   (gtwiz_init_done),
  .retry_ctr_out   (gtwiz_init_retry_ctr)
);


wire gtwiz_userclk_tx_srcclk;
wire gtwiz_userclk_tx_usrclk;
wire gtwiz_userclk_tx_usrclk2;
wire gtwiz_userclk_tx_active;
wire gtwiz_userclk_rx_srcclk;
wire gtwiz_userclk_rx_usrclk;
wire gtwiz_userclk_rx_usrclk2;
wire gtwiz_userclk_rx_active;
wire gtwiz_reset_tx_pll_and_datapath;
wire gtwiz_reset_tx_datapath;
wire gtwiz_reset_rx_pll_and_datapath = 1'b0;
wire gtwiz_reset_rx_datapath;
wire gtwiz_reset_rx_cdr_stable;
wire gtwiz_reset_tx_done;
wire gtwiz_reset_rx_done;
wire [31:0] gtwiz_userdata_tx;
wire [31:0] gtwiz_userdata_rx;
wire gtrefclk00;
wire qpll0outclk;
wire qpll0outrefclk;
wire rx8b10ben = 1'b1;
wire [0:0] rxcommadeten = 1'b1;
wire [0:0] rxmcommaalignen = 1'b1;
wire [0:0] rxpcommaalignen = 1'b1;
wire [0:0] tx8b10ben = 1'b1;
wire [15:0] txctrl0;
wire [15:0] txctrl1;
wire [7:0] txctrl2;
wire gtpowergood;
wire rxbyteisaligned;
wire rxbyterealign;
wire rxcommadet;
wire [15:0] rxctrl0;
wire [15:0] rxctrl1;
wire [7:0] rxctrl2;
wire [7:0] rxctrl3;
wire rxpmaresetdone;
wire txpmaresetdone;
wire rxrecclkout;


gty_sfp_wrapper wrapper_inst (
  .gtyrxn_in                               (gtyrxn)
 ,.gtyrxp_in                               (gtyrxp)
 ,.gtytxn_out                              (gtytxn)
 ,.gtytxp_out                              (gtytxp)
 ,.gtwiz_userclk_tx_reset_in               (gtwiz_userclk_tx_reset)
 ,.gtwiz_userclk_tx_srcclk_out             (gtwiz_userclk_tx_srcclk)
 ,.gtwiz_userclk_tx_usrclk_out             (gtwiz_userclk_tx_usrclk)
 ,.gtwiz_userclk_tx_usrclk2_out            (gtwiz_userclk_tx_usrclk2)
 ,.gtwiz_userclk_tx_active_out             (gtwiz_userclk_tx_active)
 ,.gtwiz_userclk_rx_reset_in               (gtwiz_userclk_rx_reset)
 ,.gtwiz_userclk_rx_srcclk_out             (gtwiz_userclk_rx_srcclk)
 ,.gtwiz_userclk_rx_usrclk_out             (gtwiz_userclk_rx_usrclk)
 ,.gtwiz_userclk_rx_usrclk2_out            (gtwiz_userclk_rx_usrclk2)
 ,.gtwiz_userclk_rx_active_out             (gtwiz_userclk_rx_active)
 ,.gtwiz_reset_clk_freerun_in              (gtwiz_reset_clk_freerun_buf)
 ,.gtwiz_reset_all_in                      (gtwiz_reset_all)
 ,.gtwiz_reset_tx_pll_and_datapath_in      (gtwiz_reset_tx_pll_and_datapath)
 ,.gtwiz_reset_tx_datapath_in              (gtwiz_reset_tx_datapath)
 ,.gtwiz_reset_rx_pll_and_datapath_in      (gtwiz_reset_rx_pll_and_datapath)
 ,.gtwiz_reset_rx_datapath_in              (gtwiz_reset_rx_datapath)
 ,.gtwiz_reset_rx_cdr_stable_out           (gtwiz_reset_rx_cdr_stable)
 ,.gtwiz_reset_tx_done_out                 (gtwiz_reset_tx_done)
 ,.gtwiz_reset_rx_done_out                 (gtwiz_reset_rx_done)
 ,.gtwiz_userdata_tx_in                    (gtwiz_userdata_tx)
 ,.gtwiz_userdata_rx_out                   (gtwiz_userdata_rx)
 ,.gtrefclk00_in                           (gtrefclk00)
 ,.qpll0outclk_out                         (qpll0outclk)
 ,.qpll0outrefclk_out                      (qpll0outrefclk)
 ,.rx8b10ben_in                            (rx8b10ben)
 ,.rxcommadeten_in                         (rxcommadeten)
 ,.rxmcommaalignen_in                      (rxmcommaalignen)
 ,.rxpcommaalignen_in                      (rxpcommaalignen)
 ,.tx8b10ben_in                            (tx8b10ben)
 ,.txctrl0_in                              (txctrl0)
 ,.txctrl1_in                              (txctrl1)
 ,.txctrl2_in                              (txctrl2)
 ,.gtpowergood_out                         (gtpowergood)
 ,.rxbyteisaligned_out                     (rxbyteisaligned)
 ,.rxbyterealign_out                       (rxbyterealign)
 ,.rxcommadet_out                          (rxcommadet)
 ,.rxctrl0_out                             (rxctrl0)
 ,.rxctrl1_out                             (rxctrl1)
 ,.rxctrl2_out                             (rxctrl2)
 ,.rxctrl3_out                             (rxctrl3)
 ,.rxpmaresetdone_out                      (rxpmaresetdone)
 ,.rxrecclkout_out                         (rxrecclkout)
 ,.txpmaresetdone_out                      (txpmaresetdone)
);


endmodule
