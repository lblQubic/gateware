input  DAC00_M_AXIS_ACLK
    ,input  DAC00_M_AXIS_ARESETN
    ,input  DAC00_M_AXIS_TREADY
    ,output  DAC00_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC00_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC00_M_AXIS_TSTRB
    ,output  DAC00_M_AXIS_TLAST
,input clk_dac0
,input  DAC01_M_AXIS_ACLK
    ,input  DAC01_M_AXIS_ARESETN
    ,input  DAC01_M_AXIS_TREADY
    ,output  DAC01_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC01_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC01_M_AXIS_TSTRB
    ,output  DAC01_M_AXIS_TLAST
,input  DAC02_M_AXIS_ACLK
    ,input  DAC02_M_AXIS_ARESETN
    ,input  DAC02_M_AXIS_TREADY
    ,output  DAC02_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC02_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC02_M_AXIS_TSTRB
    ,output  DAC02_M_AXIS_TLAST
,input  DAC03_M_AXIS_ACLK
    ,input  DAC03_M_AXIS_ARESETN
    ,input  DAC03_M_AXIS_TREADY
    ,output  DAC03_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC03_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC03_M_AXIS_TSTRB
    ,output  DAC03_M_AXIS_TLAST
,input  DAC10_M_AXIS_ACLK
    ,input  DAC10_M_AXIS_ARESETN
    ,input  DAC10_M_AXIS_TREADY
    ,output  DAC10_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC10_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC10_M_AXIS_TSTRB
    ,output  DAC10_M_AXIS_TLAST
,input clk_dac1
,input  DAC11_M_AXIS_ACLK
    ,input  DAC11_M_AXIS_ARESETN
    ,input  DAC11_M_AXIS_TREADY
    ,output  DAC11_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC11_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC11_M_AXIS_TSTRB
    ,output  DAC11_M_AXIS_TLAST
,input  DAC12_M_AXIS_ACLK
    ,input  DAC12_M_AXIS_ARESETN
    ,input  DAC12_M_AXIS_TREADY
    ,output  DAC12_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC12_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC12_M_AXIS_TSTRB
    ,output  DAC12_M_AXIS_TLAST
,input  DAC13_M_AXIS_ACLK
    ,input  DAC13_M_AXIS_ARESETN
    ,input  DAC13_M_AXIS_TREADY
    ,output  DAC13_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC13_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC13_M_AXIS_TSTRB
    ,output  DAC13_M_AXIS_TLAST
,input  DAC20_M_AXIS_ACLK
    ,input  DAC20_M_AXIS_ARESETN
    ,input  DAC20_M_AXIS_TREADY
    ,output  DAC20_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC20_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC20_M_AXIS_TSTRB
    ,output  DAC20_M_AXIS_TLAST
,input clk_dac2
,input  DAC21_M_AXIS_ACLK
    ,input  DAC21_M_AXIS_ARESETN
    ,input  DAC21_M_AXIS_TREADY
    ,output  DAC21_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC21_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC21_M_AXIS_TSTRB
    ,output  DAC21_M_AXIS_TLAST
,input  DAC22_M_AXIS_ACLK
    ,input  DAC22_M_AXIS_ARESETN
    ,input  DAC22_M_AXIS_TREADY
    ,output  DAC22_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC22_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC22_M_AXIS_TSTRB
    ,output  DAC22_M_AXIS_TLAST
,input  DAC23_M_AXIS_ACLK
    ,input  DAC23_M_AXIS_ARESETN
    ,input  DAC23_M_AXIS_TREADY
    ,output  DAC23_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC23_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC23_M_AXIS_TSTRB
    ,output  DAC23_M_AXIS_TLAST
,input  DAC30_M_AXIS_ACLK
    ,input  DAC30_M_AXIS_ARESETN
    ,input  DAC30_M_AXIS_TREADY
    ,output  DAC30_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC30_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC30_M_AXIS_TSTRB
    ,output  DAC30_M_AXIS_TLAST
,input clk_dac3
,input  DAC31_M_AXIS_ACLK
    ,input  DAC31_M_AXIS_ARESETN
    ,input  DAC31_M_AXIS_TREADY
    ,output  DAC31_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC31_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC31_M_AXIS_TSTRB
    ,output  DAC31_M_AXIS_TLAST
,input  DAC32_M_AXIS_ACLK
    ,input  DAC32_M_AXIS_ARESETN
    ,input  DAC32_M_AXIS_TREADY
    ,output  DAC32_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC32_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC32_M_AXIS_TSTRB
    ,output  DAC32_M_AXIS_TLAST
,input  DAC33_M_AXIS_ACLK
    ,input  DAC33_M_AXIS_ARESETN
    ,input  DAC33_M_AXIS_TREADY
    ,output  DAC33_M_AXIS_TVALID
    ,output  [DAC_AXIS_DATAWIDTH-1 : 0] DAC33_M_AXIS_TDATA
    ,output  [(DAC_AXIS_DATAWIDTH/8)-1 : 0] DAC33_M_AXIS_TSTRB
    ,output  DAC33_M_AXIS_TLAST
,input  ADC00_S_AXIS_ACLK
    ,input  ADC00_S_AXIS_ARESETN
    ,output  ADC00_S_AXIS_TREADY
    ,input  ADC00_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC00_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC00_S_AXIS_TSTRB
    ,input  ADC00_S_AXIS_TLAST
,input clk_adc0
,input  ADC01_S_AXIS_ACLK
    ,input  ADC01_S_AXIS_ARESETN
    ,output  ADC01_S_AXIS_TREADY
    ,input  ADC01_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC01_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC01_S_AXIS_TSTRB
    ,input  ADC01_S_AXIS_TLAST
,input  ADC02_S_AXIS_ACLK
    ,input  ADC02_S_AXIS_ARESETN
    ,output  ADC02_S_AXIS_TREADY
    ,input  ADC02_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC02_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC02_S_AXIS_TSTRB
    ,input  ADC02_S_AXIS_TLAST
,input  ADC03_S_AXIS_ACLK
    ,input  ADC03_S_AXIS_ARESETN
    ,output  ADC03_S_AXIS_TREADY
    ,input  ADC03_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC03_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC03_S_AXIS_TSTRB
    ,input  ADC03_S_AXIS_TLAST
,input  ADC10_S_AXIS_ACLK
    ,input  ADC10_S_AXIS_ARESETN
    ,output  ADC10_S_AXIS_TREADY
    ,input  ADC10_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC10_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC10_S_AXIS_TSTRB
    ,input  ADC10_S_AXIS_TLAST
,input clk_adc1
,input  ADC11_S_AXIS_ACLK
    ,input  ADC11_S_AXIS_ARESETN
    ,output  ADC11_S_AXIS_TREADY
    ,input  ADC11_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC11_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC11_S_AXIS_TSTRB
    ,input  ADC11_S_AXIS_TLAST
,input  ADC12_S_AXIS_ACLK
    ,input  ADC12_S_AXIS_ARESETN
    ,output  ADC12_S_AXIS_TREADY
    ,input  ADC12_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC12_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC12_S_AXIS_TSTRB
    ,input  ADC12_S_AXIS_TLAST
,input  ADC13_S_AXIS_ACLK
    ,input  ADC13_S_AXIS_ARESETN
    ,output  ADC13_S_AXIS_TREADY
    ,input  ADC13_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC13_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC13_S_AXIS_TSTRB
    ,input  ADC13_S_AXIS_TLAST
,input  ADC20_S_AXIS_ACLK
    ,input  ADC20_S_AXIS_ARESETN
    ,output  ADC20_S_AXIS_TREADY
    ,input  ADC20_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC20_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC20_S_AXIS_TSTRB
    ,input  ADC20_S_AXIS_TLAST
,input clk_adc2
,input  ADC21_S_AXIS_ACLK
    ,input  ADC21_S_AXIS_ARESETN
    ,output  ADC21_S_AXIS_TREADY
    ,input  ADC21_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC21_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC21_S_AXIS_TSTRB
    ,input  ADC21_S_AXIS_TLAST
,input  ADC22_S_AXIS_ACLK
    ,input  ADC22_S_AXIS_ARESETN
    ,output  ADC22_S_AXIS_TREADY
    ,input  ADC22_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC22_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC22_S_AXIS_TSTRB
    ,input  ADC22_S_AXIS_TLAST
,input  ADC23_S_AXIS_ACLK
    ,input  ADC23_S_AXIS_ARESETN
    ,output  ADC23_S_AXIS_TREADY
    ,input  ADC23_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC23_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC23_S_AXIS_TSTRB
    ,input  ADC23_S_AXIS_TLAST
,input  ADC30_S_AXIS_ACLK
    ,input  ADC30_S_AXIS_ARESETN
    ,output  ADC30_S_AXIS_TREADY
    ,input  ADC30_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC30_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC30_S_AXIS_TSTRB
    ,input  ADC30_S_AXIS_TLAST
,input clk_adc3
,input  ADC31_S_AXIS_ACLK
    ,input  ADC31_S_AXIS_ARESETN
    ,output  ADC31_S_AXIS_TREADY
    ,input  ADC31_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC31_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC31_S_AXIS_TSTRB
    ,input  ADC31_S_AXIS_TLAST
,input  ADC32_S_AXIS_ACLK
    ,input  ADC32_S_AXIS_ARESETN
    ,output  ADC32_S_AXIS_TREADY
    ,input  ADC32_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC32_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC32_S_AXIS_TSTRB
    ,input  ADC32_S_AXIS_TLAST
,input  ADC33_S_AXIS_ACLK
    ,input  ADC33_S_AXIS_ARESETN
    ,output  ADC33_S_AXIS_TREADY
    ,input  ADC33_S_AXIS_TVALID
    ,input  [ADC_AXIS_DATAWIDTH-1 : 0] ADC33_S_AXIS_TDATA
    ,input  [(ADC_AXIS_DATAWIDTH/8)-1 : 0] ADC33_S_AXIS_TSTRB
    ,input  ADC33_S_AXIS_TLAST