.LB1_DATAWIDTH(LB1_DATAWIDTH),.LB1_ADDRWIDTH(LB1_ADDRWIDTH)
,.LB2_DATAWIDTH(LB2_DATAWIDTH),.LB2_ADDRWIDTH(LB2_ADDRWIDTH)
,.LB3_DATAWIDTH(LB3_DATAWIDTH),.LB3_ADDRWIDTH(LB3_ADDRWIDTH)
,.LB4_DATAWIDTH(LB4_DATAWIDTH),.LB4_ADDRWIDTH(LB4_ADDRWIDTH)
,.DAC_AXIS_DATAWIDTH(DAC_AXIS_DATAWIDTH)
,`include "bram_parainst.vh"
