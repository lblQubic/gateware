module ilaauto (input clk
,input [32-1:0] probe0
,input [16-1:0] probe1
,input [1-1:0] probe2
);
endmodule
