parameter INIT_acqbuf0=""
,parameter INIT_acqbuf1=""
,parameter INIT_command0=""
,parameter INIT_command1=""
,parameter INIT_command2=""
,parameter INIT_qdrvfreq0=""
,parameter INIT_qdrvfreq1=""
,parameter INIT_qdrvfreq2=""
,parameter INIT_rdrvfreq0=""
,parameter INIT_rdrvfreq1=""
,parameter INIT_rdrvfreq2=""
,parameter INIT_dacmon0=""
,parameter INIT_dacmon1=""
,parameter INIT_dacmon2=""
,parameter INIT_dacmon3=""
,parameter INIT_qdrvenv0=""
,parameter INIT_qdrvenv1=""
,parameter INIT_qdrvenv2=""
,parameter INIT_rdloenv0=""
,parameter INIT_rdloenv1=""
,parameter INIT_rdloenv2=""
,parameter INIT_rdrvenv0=""
,parameter INIT_rdrvenv1=""
,parameter INIT_rdrvenv2=""
,parameter INIT_accbuf0=""
,parameter INIT_accbuf1=""
,parameter INIT_accbuf2=""
,parameter INIT_rdlofreq0=""
,parameter INIT_rdlofreq1=""
,parameter INIT_rdlofreq2=""