module ilaauto (input clk
,input [32-1:0] probe0
,input [1-1:0] probe1
,input [1-1:0] probe2
,input [256-1:0] probe3
,input [32-1:0] probe4
,input [1-1:0] probe5
,input [1-1:0] probe6
,input [256-1:0] probe7
);
endmodule
