.acqbuf0_W(acqbuf0_W)
,.acqbuf1_W(acqbuf1_W)
,.command0_R(command0_R)
,.command1_R(command1_R)
,.command2_R(command2_R)
,.command3_R(command3_R)
,.command4_R(command4_R)
,.command5_R(command5_R)
,.command6_R(command6_R)
,.command7_R(command7_R)
,.qdrvfreq0_R(qdrvfreq0_R)
,.qdrvfreq1_R(qdrvfreq1_R)
,.qdrvfreq2_R(qdrvfreq2_R)
,.qdrvfreq3_R(qdrvfreq3_R)
,.qdrvfreq4_R(qdrvfreq4_R)
,.qdrvfreq5_R(qdrvfreq5_R)
,.qdrvfreq6_R(qdrvfreq6_R)
,.qdrvfreq7_R(qdrvfreq7_R)
,.rdrvfreq0_R(rdrvfreq0_R)
,.rdrvfreq1_R(rdrvfreq1_R)
,.rdrvfreq2_R(rdrvfreq2_R)
,.rdrvfreq3_R(rdrvfreq3_R)
,.rdrvfreq4_R(rdrvfreq4_R)
,.rdrvfreq5_R(rdrvfreq5_R)
,.rdrvfreq6_R(rdrvfreq6_R)
,.rdrvfreq7_R(rdrvfreq7_R)
,.dacmon0_W(dacmon0_W)
,.dacmon1_W(dacmon1_W)
,.dacmon2_W(dacmon2_W)
,.dacmon3_W(dacmon3_W)
,.qdrvenv0_R(qdrvenv0_R)
,.qdrvenv1_R(qdrvenv1_R)
,.qdrvenv2_R(qdrvenv2_R)
,.qdrvenv3_R(qdrvenv3_R)
,.qdrvenv4_R(qdrvenv4_R)
,.qdrvenv5_R(qdrvenv5_R)
,.qdrvenv6_R(qdrvenv6_R)
,.qdrvenv7_R(qdrvenv7_R)
,.rdloenv0_R(rdloenv0_R)
,.rdloenv1_R(rdloenv1_R)
,.rdloenv2_R(rdloenv2_R)
,.rdloenv3_R(rdloenv3_R)
,.rdloenv4_R(rdloenv4_R)
,.rdloenv5_R(rdloenv5_R)
,.rdloenv6_R(rdloenv6_R)
,.rdloenv7_R(rdloenv7_R)
,.rdrvenv0_R(rdrvenv0_R)
,.rdrvenv1_R(rdrvenv1_R)
,.rdrvenv2_R(rdrvenv2_R)
,.rdrvenv3_R(rdrvenv3_R)
,.rdrvenv4_R(rdrvenv4_R)
,.rdrvenv5_R(rdrvenv5_R)
,.rdrvenv6_R(rdrvenv6_R)
,.rdrvenv7_R(rdrvenv7_R)
,.accbuf0_W(accbuf0_W)
,.accbuf1_W(accbuf1_W)
,.accbuf2_W(accbuf2_W)
,.accbuf3_W(accbuf3_W)
,.accbuf4_W(accbuf4_W)
,.accbuf5_W(accbuf5_W)
,.accbuf6_W(accbuf6_W)
,.accbuf7_W(accbuf7_W)
,.rdlofreq0_R(rdlofreq0_R)
,.rdlofreq1_R(rdlofreq1_R)
,.rdlofreq2_R(rdlofreq2_R)
,.rdlofreq3_R(rdlofreq3_R)
,.rdlofreq4_R(rdlofreq4_R)
,.rdlofreq5_R(rdlofreq5_R)
,.rdlofreq6_R(rdlofreq6_R)
,.rdlofreq7_R(rdlofreq7_R)
,.sdbuf0_W(sdbuf0_W)
,.sdbuf1_W(sdbuf1_W)
,.sdbuf2_W(sdbuf2_W)
,.sdbuf3_W(sdbuf3_W)
,.sdbuf4_W(sdbuf4_W)
,.sdbuf5_W(sdbuf5_W)
,.sdbuf6_W(sdbuf6_W)
,.sdbuf7_W(sdbuf7_W)