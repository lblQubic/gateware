.acqbuf0_R(acqbuf0_R)
,.acqbuf1_R(acqbuf1_R)
,.command0_W(command0_W)
,.command1_W(command1_W)
,.command2_W(command2_W)
,.qdrvfreq0_W(qdrvfreq0_W)
,.qdrvfreq1_W(qdrvfreq1_W)
,.qdrvfreq2_W(qdrvfreq2_W)
,.rdrvfreq0_W(rdrvfreq0_W)
,.rdrvfreq1_W(rdrvfreq1_W)
,.rdrvfreq2_W(rdrvfreq2_W)
,.dacmon0_R(dacmon0_R)
,.dacmon1_R(dacmon1_R)
,.dacmon2_R(dacmon2_R)
,.dacmon3_R(dacmon3_R)
,.qdrvenv0_W(qdrvenv0_W)
,.qdrvenv1_W(qdrvenv1_W)
,.qdrvenv2_W(qdrvenv2_W)
,.rdloenv0_W(rdloenv0_W)
,.rdloenv1_W(rdloenv1_W)
,.rdloenv2_W(rdloenv2_W)
,.rdrvenv0_W(rdrvenv0_W)
,.rdrvenv1_W(rdrvenv1_W)
,.rdrvenv2_W(rdrvenv2_W)
,.accbuf0_R(accbuf0_R)
,.accbuf1_R(accbuf1_R)
,.accbuf2_R(accbuf2_R)
,.rdlofreq0_W(rdlofreq0_W)
,.rdlofreq1_W(rdlofreq1_W)
,.rdlofreq2_W(rdlofreq2_W)