ifbram acqbuf0_R
,ifbram acqbuf1_R
,ifbram command0_W
,ifbram command1_W
,ifbram command2_W
,ifbram qdrvfreq0_W
,ifbram qdrvfreq1_W
,ifbram qdrvfreq2_W
,ifbram rdrvfreq0_W
,ifbram rdrvfreq1_W
,ifbram rdrvfreq2_W
,ifbram dacmon0_R
,ifbram dacmon1_R
,ifbram dacmon2_R
,ifbram dacmon3_R
,ifbram qdrvenv0_W
,ifbram qdrvenv1_W
,ifbram qdrvenv2_W
,ifbram rdloenv0_W
,ifbram rdloenv1_W
,ifbram rdloenv2_W
,ifbram rdrvenv0_W
,ifbram rdrvenv1_W
,ifbram rdrvenv2_W
,ifbram accbuf0_R
,ifbram accbuf1_R
,ifbram accbuf2_R
,ifbram rdlofreq0_W
,ifbram rdlofreq1_W
,ifbram rdlofreq2_W