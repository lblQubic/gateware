ifbram acqbuf0_W
,ifbram acqbuf1_W
,ifbram command0_R
,ifbram command1_R
,ifbram command2_R
,ifbram qdrvfreq0_R
,ifbram qdrvfreq1_R
,ifbram qdrvfreq2_R
,ifbram rdrvfreq0_R
,ifbram rdrvfreq1_R
,ifbram rdrvfreq2_R
,ifbram dacmon0_W
,ifbram dacmon1_W
,ifbram dacmon2_W
,ifbram dacmon3_W
,ifbram qdrvenv0_R
,ifbram qdrvenv1_R
,ifbram qdrvenv2_R
,ifbram rdloenv0_R
,ifbram rdloenv1_R
,ifbram rdloenv2_R
,ifbram rdrvenv0_R
,ifbram rdrvenv1_R
,ifbram rdrvenv2_R
,ifbram accbuf0_W
,ifbram accbuf1_W
,ifbram accbuf2_W
,ifbram rdlofreq0_R
,ifbram rdlofreq1_R
,ifbram rdlofreq2_R