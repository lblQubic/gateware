output ACCBUF0_clk
,output ACCBUF0_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF0_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF0_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF0_dout
,output ACCBUF0_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF0_we

,output ACCBUF1_clk
,output ACCBUF1_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF1_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF1_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF1_dout
,output ACCBUF1_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF1_we

,output ACCBUF2_clk
,output ACCBUF2_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF2_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF2_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF2_dout
,output ACCBUF2_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF2_we

,output ACCBUF3_clk
,output ACCBUF3_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF3_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF3_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF3_dout
,output ACCBUF3_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF3_we

,output ACCBUF4_clk
,output ACCBUF4_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF4_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF4_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF4_dout
,output ACCBUF4_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF4_we

,output ACCBUF5_clk
,output ACCBUF5_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF5_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF5_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF5_dout
,output ACCBUF5_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF5_we

,output ACCBUF6_clk
,output ACCBUF6_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF6_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF6_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF6_dout
,output ACCBUF6_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF6_we

,output ACCBUF7_clk
,output ACCBUF7_rst
,output [BRAMADDRWIDTH-1:0] ACCBUF7_addr
,output [ACCBUF_DATAWIDTH-1:0] ACCBUF7_din
,input [ACCBUF_DATAWIDTH-1:0] ACCBUF7_dout
,output ACCBUF7_en
,output [ACCBUF_DATAWIDTH/8-1:0] ACCBUF7_we

,output ACQBUF0_clk
,output ACQBUF0_rst
,output [BRAMADDRWIDTH-1:0] ACQBUF0_addr
,output [ACQBUF_DATAWIDTH-1:0] ACQBUF0_din
,input [ACQBUF_DATAWIDTH-1:0] ACQBUF0_dout
,output ACQBUF0_en
,output [ACQBUF_DATAWIDTH/8-1:0] ACQBUF0_we

,output ACQBUF1_clk
,output ACQBUF1_rst
,output [BRAMADDRWIDTH-1:0] ACQBUF1_addr
,output [ACQBUF_DATAWIDTH-1:0] ACQBUF1_din
,input [ACQBUF_DATAWIDTH-1:0] ACQBUF1_dout
,output ACQBUF1_en
,output [ACQBUF_DATAWIDTH/8-1:0] ACQBUF1_we

,output COMMAND0_clk
,output COMMAND0_rst
,output [BRAMADDRWIDTH-1:0] COMMAND0_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND0_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND0_dout
,output COMMAND0_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND0_we

,output COMMAND1_clk
,output COMMAND1_rst
,output [BRAMADDRWIDTH-1:0] COMMAND1_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND1_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND1_dout
,output COMMAND1_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND1_we

,output COMMAND2_clk
,output COMMAND2_rst
,output [BRAMADDRWIDTH-1:0] COMMAND2_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND2_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND2_dout
,output COMMAND2_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND2_we

,output COMMAND3_clk
,output COMMAND3_rst
,output [BRAMADDRWIDTH-1:0] COMMAND3_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND3_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND3_dout
,output COMMAND3_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND3_we

,output COMMAND4_clk
,output COMMAND4_rst
,output [BRAMADDRWIDTH-1:0] COMMAND4_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND4_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND4_dout
,output COMMAND4_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND4_we

,output COMMAND5_clk
,output COMMAND5_rst
,output [BRAMADDRWIDTH-1:0] COMMAND5_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND5_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND5_dout
,output COMMAND5_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND5_we

,output COMMAND6_clk
,output COMMAND6_rst
,output [BRAMADDRWIDTH-1:0] COMMAND6_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND6_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND6_dout
,output COMMAND6_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND6_we

,output COMMAND7_clk
,output COMMAND7_rst
,output [BRAMADDRWIDTH-1:0] COMMAND7_addr
,output [COMMAND_DATAWIDTH-1:0] COMMAND7_din
,input [COMMAND_DATAWIDTH-1:0] COMMAND7_dout
,output COMMAND7_en
,output [COMMAND_DATAWIDTH/8-1:0] COMMAND7_we

,output DACMON0_clk
,output DACMON0_rst
,output [BRAMADDRWIDTH-1:0] DACMON0_addr
,output [DACMON_DATAWIDTH-1:0] DACMON0_din
,input [DACMON_DATAWIDTH-1:0] DACMON0_dout
,output DACMON0_en
,output [DACMON_DATAWIDTH/8-1:0] DACMON0_we

,output DACMON1_clk
,output DACMON1_rst
,output [BRAMADDRWIDTH-1:0] DACMON1_addr
,output [DACMON_DATAWIDTH-1:0] DACMON1_din
,input [DACMON_DATAWIDTH-1:0] DACMON1_dout
,output DACMON1_en
,output [DACMON_DATAWIDTH/8-1:0] DACMON1_we

,output DACMON2_clk
,output DACMON2_rst
,output [BRAMADDRWIDTH-1:0] DACMON2_addr
,output [DACMON_DATAWIDTH-1:0] DACMON2_din
,input [DACMON_DATAWIDTH-1:0] DACMON2_dout
,output DACMON2_en
,output [DACMON_DATAWIDTH/8-1:0] DACMON2_we

,output DACMON3_clk
,output DACMON3_rst
,output [BRAMADDRWIDTH-1:0] DACMON3_addr
,output [DACMON_DATAWIDTH-1:0] DACMON3_din
,input [DACMON_DATAWIDTH-1:0] DACMON3_dout
,output DACMON3_en
,output [DACMON_DATAWIDTH/8-1:0] DACMON3_we

,output QDRVENV0_clk
,output QDRVENV0_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV0_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV0_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV0_dout
,output QDRVENV0_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV0_we

,output QDRVENV1_clk
,output QDRVENV1_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV1_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV1_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV1_dout
,output QDRVENV1_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV1_we

,output QDRVENV2_clk
,output QDRVENV2_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV2_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV2_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV2_dout
,output QDRVENV2_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV2_we

,output QDRVENV3_clk
,output QDRVENV3_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV3_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV3_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV3_dout
,output QDRVENV3_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV3_we

,output QDRVENV4_clk
,output QDRVENV4_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV4_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV4_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV4_dout
,output QDRVENV4_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV4_we

,output QDRVENV5_clk
,output QDRVENV5_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV5_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV5_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV5_dout
,output QDRVENV5_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV5_we

,output QDRVENV6_clk
,output QDRVENV6_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV6_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV6_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV6_dout
,output QDRVENV6_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV6_we

,output QDRVENV7_clk
,output QDRVENV7_rst
,output [BRAMADDRWIDTH-1:0] QDRVENV7_addr
,output [QDRVENV_DATAWIDTH-1:0] QDRVENV7_din
,input [QDRVENV_DATAWIDTH-1:0] QDRVENV7_dout
,output QDRVENV7_en
,output [QDRVENV_DATAWIDTH/8-1:0] QDRVENV7_we

,output QDRVFREQ0_clk
,output QDRVFREQ0_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ0_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ0_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ0_dout
,output QDRVFREQ0_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ0_we

,output QDRVFREQ1_clk
,output QDRVFREQ1_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ1_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ1_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ1_dout
,output QDRVFREQ1_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ1_we

,output QDRVFREQ2_clk
,output QDRVFREQ2_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ2_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ2_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ2_dout
,output QDRVFREQ2_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ2_we

,output QDRVFREQ3_clk
,output QDRVFREQ3_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ3_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ3_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ3_dout
,output QDRVFREQ3_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ3_we

,output QDRVFREQ4_clk
,output QDRVFREQ4_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ4_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ4_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ4_dout
,output QDRVFREQ4_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ4_we

,output QDRVFREQ5_clk
,output QDRVFREQ5_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ5_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ5_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ5_dout
,output QDRVFREQ5_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ5_we

,output QDRVFREQ6_clk
,output QDRVFREQ6_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ6_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ6_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ6_dout
,output QDRVFREQ6_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ6_we

,output QDRVFREQ7_clk
,output QDRVFREQ7_rst
,output [BRAMADDRWIDTH-1:0] QDRVFREQ7_addr
,output [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ7_din
,input [QDRVFREQ_DATAWIDTH-1:0] QDRVFREQ7_dout
,output QDRVFREQ7_en
,output [QDRVFREQ_DATAWIDTH/8-1:0] QDRVFREQ7_we

,output RDLOENV0_clk
,output RDLOENV0_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV0_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV0_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV0_dout
,output RDLOENV0_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV0_we

,output RDLOENV1_clk
,output RDLOENV1_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV1_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV1_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV1_dout
,output RDLOENV1_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV1_we

,output RDLOENV2_clk
,output RDLOENV2_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV2_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV2_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV2_dout
,output RDLOENV2_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV2_we

,output RDLOENV3_clk
,output RDLOENV3_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV3_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV3_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV3_dout
,output RDLOENV3_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV3_we

,output RDLOENV4_clk
,output RDLOENV4_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV4_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV4_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV4_dout
,output RDLOENV4_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV4_we

,output RDLOENV5_clk
,output RDLOENV5_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV5_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV5_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV5_dout
,output RDLOENV5_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV5_we

,output RDLOENV6_clk
,output RDLOENV6_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV6_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV6_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV6_dout
,output RDLOENV6_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV6_we

,output RDLOENV7_clk
,output RDLOENV7_rst
,output [BRAMADDRWIDTH-1:0] RDLOENV7_addr
,output [RDLOENV_DATAWIDTH-1:0] RDLOENV7_din
,input [RDLOENV_DATAWIDTH-1:0] RDLOENV7_dout
,output RDLOENV7_en
,output [RDLOENV_DATAWIDTH/8-1:0] RDLOENV7_we

,output RDLOFREQ0_clk
,output RDLOFREQ0_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ0_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ0_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ0_dout
,output RDLOFREQ0_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ0_we

,output RDLOFREQ1_clk
,output RDLOFREQ1_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ1_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ1_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ1_dout
,output RDLOFREQ1_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ1_we

,output RDLOFREQ2_clk
,output RDLOFREQ2_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ2_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ2_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ2_dout
,output RDLOFREQ2_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ2_we

,output RDLOFREQ3_clk
,output RDLOFREQ3_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ3_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ3_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ3_dout
,output RDLOFREQ3_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ3_we

,output RDLOFREQ4_clk
,output RDLOFREQ4_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ4_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ4_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ4_dout
,output RDLOFREQ4_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ4_we

,output RDLOFREQ5_clk
,output RDLOFREQ5_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ5_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ5_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ5_dout
,output RDLOFREQ5_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ5_we

,output RDLOFREQ6_clk
,output RDLOFREQ6_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ6_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ6_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ6_dout
,output RDLOFREQ6_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ6_we

,output RDLOFREQ7_clk
,output RDLOFREQ7_rst
,output [BRAMADDRWIDTH-1:0] RDLOFREQ7_addr
,output [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ7_din
,input [RDLOFREQ_DATAWIDTH-1:0] RDLOFREQ7_dout
,output RDLOFREQ7_en
,output [RDLOFREQ_DATAWIDTH/8-1:0] RDLOFREQ7_we

,output RDRVENV0_clk
,output RDRVENV0_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV0_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV0_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV0_dout
,output RDRVENV0_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV0_we

,output RDRVENV1_clk
,output RDRVENV1_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV1_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV1_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV1_dout
,output RDRVENV1_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV1_we

,output RDRVENV2_clk
,output RDRVENV2_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV2_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV2_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV2_dout
,output RDRVENV2_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV2_we

,output RDRVENV3_clk
,output RDRVENV3_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV3_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV3_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV3_dout
,output RDRVENV3_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV3_we

,output RDRVENV4_clk
,output RDRVENV4_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV4_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV4_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV4_dout
,output RDRVENV4_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV4_we

,output RDRVENV5_clk
,output RDRVENV5_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV5_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV5_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV5_dout
,output RDRVENV5_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV5_we

,output RDRVENV6_clk
,output RDRVENV6_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV6_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV6_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV6_dout
,output RDRVENV6_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV6_we

,output RDRVENV7_clk
,output RDRVENV7_rst
,output [BRAMADDRWIDTH-1:0] RDRVENV7_addr
,output [RDRVENV_DATAWIDTH-1:0] RDRVENV7_din
,input [RDRVENV_DATAWIDTH-1:0] RDRVENV7_dout
,output RDRVENV7_en
,output [RDRVENV_DATAWIDTH/8-1:0] RDRVENV7_we

,output RDRVFREQ0_clk
,output RDRVFREQ0_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ0_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ0_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ0_dout
,output RDRVFREQ0_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ0_we

,output RDRVFREQ1_clk
,output RDRVFREQ1_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ1_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ1_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ1_dout
,output RDRVFREQ1_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ1_we

,output RDRVFREQ2_clk
,output RDRVFREQ2_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ2_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ2_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ2_dout
,output RDRVFREQ2_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ2_we

,output RDRVFREQ3_clk
,output RDRVFREQ3_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ3_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ3_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ3_dout
,output RDRVFREQ3_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ3_we

,output RDRVFREQ4_clk
,output RDRVFREQ4_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ4_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ4_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ4_dout
,output RDRVFREQ4_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ4_we

,output RDRVFREQ5_clk
,output RDRVFREQ5_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ5_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ5_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ5_dout
,output RDRVFREQ5_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ5_we

,output RDRVFREQ6_clk
,output RDRVFREQ6_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ6_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ6_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ6_dout
,output RDRVFREQ6_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ6_we

,output RDRVFREQ7_clk
,output RDRVFREQ7_rst
,output [BRAMADDRWIDTH-1:0] RDRVFREQ7_addr
,output [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ7_din
,input [RDRVFREQ_DATAWIDTH-1:0] RDRVFREQ7_dout
,output RDRVFREQ7_en
,output [RDRVFREQ_DATAWIDTH/8-1:0] RDRVFREQ7_we

,output SDBUF0_clk
,output SDBUF0_rst
,output [BRAMADDRWIDTH-1:0] SDBUF0_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF0_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF0_dout
,output SDBUF0_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF0_we

,output SDBUF1_clk
,output SDBUF1_rst
,output [BRAMADDRWIDTH-1:0] SDBUF1_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF1_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF1_dout
,output SDBUF1_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF1_we

,output SDBUF2_clk
,output SDBUF2_rst
,output [BRAMADDRWIDTH-1:0] SDBUF2_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF2_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF2_dout
,output SDBUF2_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF2_we

,output SDBUF3_clk
,output SDBUF3_rst
,output [BRAMADDRWIDTH-1:0] SDBUF3_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF3_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF3_dout
,output SDBUF3_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF3_we

,output SDBUF4_clk
,output SDBUF4_rst
,output [BRAMADDRWIDTH-1:0] SDBUF4_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF4_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF4_dout
,output SDBUF4_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF4_we

,output SDBUF5_clk
,output SDBUF5_rst
,output [BRAMADDRWIDTH-1:0] SDBUF5_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF5_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF5_dout
,output SDBUF5_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF5_we

,output SDBUF6_clk
,output SDBUF6_rst
,output [BRAMADDRWIDTH-1:0] SDBUF6_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF6_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF6_dout
,output SDBUF6_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF6_we

,output SDBUF7_clk
,output SDBUF7_rst
,output [BRAMADDRWIDTH-1:0] SDBUF7_addr
,output [SDBUF_DATAWIDTH-1:0] SDBUF7_din
,input [SDBUF_DATAWIDTH-1:0] SDBUF7_dout
,output SDBUF7_en
,output [SDBUF_DATAWIDTH/8-1:0] SDBUF7_we
