parameter NCFGRESETN=8
,parameter NDSPRESETN=42
,parameter NPSRESETN=3
,parameter NADC3RESETN=1