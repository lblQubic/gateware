.LB_DATAWIDTH(LB_DATAWIDTH)
,.LB_ADDRWIDTH(LB_ADDRWIDTH)
,.DAC_AXIS_DATAWIDTH(DAC_AXIS_DATAWIDTH)
,`include "bram_parainst.vh"
