	.aresetn( aresetn )
	,.pl_clk0( pl_clk0 )
,.cfgresetn00( cfgresetn00 )
,.cfgresetn01( cfgresetn01 )
,.cfgresetn02( cfgresetn02 )
,.cfgresetn03( cfgresetn03 )
,.cfgresetn04( cfgresetn04 )
,.cfgresetn05( cfgresetn05 )
,.cfgresetn06( cfgresetn06 )
,.cfgresetn07( cfgresetn07 )
,.cfgresetn08( cfgresetn08 )
,.cfgresetn09( cfgresetn09 )
,.cfgresetn10( cfgresetn10 )
,.cfgresetn11( cfgresetn11 )
,.cfgresetn12( cfgresetn12 )
,.cfgresetn13( cfgresetn13 )
,.cfgresetn14( cfgresetn14 )
,.cfgresetn15( cfgresetn15 )
,.cfgresetn16( cfgresetn16 )
,.cfgresetn17( cfgresetn17 )
,.cfgresetn18( cfgresetn18 )
,.cfgresetn19( cfgresetn19 )
,.cfgresetn20( cfgresetn20 )
,.cfgresetn21( cfgresetn21 )
,.cfgresetn22( cfgresetn22 )
,.cfgresetn23( cfgresetn23 )
,.cfgresetn24( cfgresetn24 )
,.cfgresetn25( cfgresetn25 )
,.cfgresetn26( cfgresetn26 )
,.cfgresetn27( cfgresetn27 )
,.cfgresetn28( cfgresetn28 )
,.cfgresetn29( cfgresetn29 )

,.dspresetn00( dspresetn00 )
,.dspresetn01( dspresetn01 )
,.dspresetn02( dspresetn02 )
,.dspresetn03( dspresetn03 )
,.dspresetn04( dspresetn04 )
,.dspresetn05( dspresetn05 )
,.dspresetn06( dspresetn06 )
,.dspresetn07( dspresetn07 )


,.psresetn00( psresetn00 )
,.psresetn01( psresetn01 )
,.psresetn02( psresetn02 )
,.adc2resetn00( adc2resetn00 )
,.adc2resetn01( adc2resetn01 )
,.adc2resetn02( adc2resetn02 )


,.lb1_wren( lb1_wren )
,.lb1_rden( lb1_rden )
,.lb1_waddr( lb1_waddr )
,.lb1_wdata( lb1_wdata )
,.lb1_raddr( lb1_raddr )
,.lb1_rdata( lb1_rdata )
,.lb1_rvalid( lb1_rvalid )
,.lb1_clk( lb1_clk )
,.lb1_aresetn( lb1_aresetn )
,.lb2_wren( lb2_wren )
,.lb2_rden( lb2_rden )
,.lb2_waddr( lb2_waddr )
,.lb2_wdata( lb2_wdata )
,.lb2_raddr( lb2_raddr )
,.lb2_rdata( lb2_rdata )
,.lb2_rvalid( lb2_rvalid )
,.lb2_clk( lb2_clk )
,.lb2_aresetn( lb2_aresetn )
,.BRAM_TOHOST0_clk( BRAM_TOHOST0_clk )
,.BRAM_TOHOST0_rst( BRAM_TOHOST0_rst )
,.BRAM_TOHOST0_addr( BRAM_TOHOST0_addr )
,.BRAM_TOHOST0_din( BRAM_TOHOST0_din )
,.BRAM_TOHOST0_dout( BRAM_TOHOST0_dout )
,.BRAM_TOHOST0_en( BRAM_TOHOST0_en )
,.BRAM_TOHOST0_we( BRAM_TOHOST0_we )
//,.bram_rsta_busy( bram_rsta_busy )
//,.bram_rstb_busy( bram_rstb_busy )
,.BRAM_TOHOST1_clk( BRAM_TOHOST1_clk )
,.BRAM_TOHOST1_rst( BRAM_TOHOST1_rst )
,.BRAM_TOHOST1_addr( BRAM_TOHOST1_addr )
,.BRAM_TOHOST1_din( BRAM_TOHOST1_din )
,.BRAM_TOHOST1_dout( BRAM_TOHOST1_dout )
,.BRAM_TOHOST1_en( BRAM_TOHOST1_en )
,.BRAM_TOHOST1_we( BRAM_TOHOST1_we )


,.BRAM_FROMHOST0_clk( BRAM_FROMHOST0_clk )
,.BRAM_FROMHOST0_rst( BRAM_FROMHOST0_rst )
,.BRAM_FROMHOST0_addr( BRAM_FROMHOST0_addr )
,.BRAM_FROMHOST0_din( BRAM_FROMHOST0_din )
,.BRAM_FROMHOST0_dout( BRAM_FROMHOST0_dout )
,.BRAM_FROMHOST0_en( BRAM_FROMHOST0_en )
,.BRAM_FROMHOST0_we( BRAM_FROMHOST0_we )
,.BRAM_FROMHOST1_clk( BRAM_FROMHOST1_clk )
,.BRAM_FROMHOST1_rst( BRAM_FROMHOST1_rst )
,.BRAM_FROMHOST1_addr( BRAM_FROMHOST1_addr )
,.BRAM_FROMHOST1_din( BRAM_FROMHOST1_din )
,.BRAM_FROMHOST1_dout( BRAM_FROMHOST1_dout )
,.BRAM_FROMHOST1_en( BRAM_FROMHOST1_en )
,.BRAM_FROMHOST1_we( BRAM_FROMHOST1_we )

,.BRAM_FROMHOST2_clk( BRAM_FROMHOST2_clk )
,.BRAM_FROMHOST2_rst( BRAM_FROMHOST2_rst )
,.BRAM_FROMHOST2_addr( BRAM_FROMHOST2_addr )
,.BRAM_FROMHOST2_din( BRAM_FROMHOST2_din )
,.BRAM_FROMHOST2_dout( BRAM_FROMHOST2_dout )
,.BRAM_FROMHOST2_en( BRAM_FROMHOST2_en )
,.BRAM_FROMHOST2_we( BRAM_FROMHOST2_we )
,.BRAM_FROMHOST3_clk( BRAM_FROMHOST3_clk )
,.BRAM_FROMHOST3_rst( BRAM_FROMHOST3_rst )
,.BRAM_FROMHOST3_addr( BRAM_FROMHOST3_addr )
,.BRAM_FROMHOST3_din( BRAM_FROMHOST3_din )
,.BRAM_FROMHOST3_dout( BRAM_FROMHOST3_dout )
,.BRAM_FROMHOST3_en( BRAM_FROMHOST3_en )
,.BRAM_FROMHOST3_we( BRAM_FROMHOST3_we )

,.BRAM_FROMHOST4_clk( BRAM_FROMHOST4_clk )
,.BRAM_FROMHOST4_rst( BRAM_FROMHOST4_rst )
,.BRAM_FROMHOST4_addr( BRAM_FROMHOST4_addr )
,.BRAM_FROMHOST4_din( BRAM_FROMHOST4_din )
,.BRAM_FROMHOST4_dout( BRAM_FROMHOST4_dout )
,.BRAM_FROMHOST4_en( BRAM_FROMHOST4_en )
,.BRAM_FROMHOST4_we( BRAM_FROMHOST4_we )

,.BRAM_FROMHOST5_clk( BRAM_FROMHOST5_clk )
,.BRAM_FROMHOST5_rst( BRAM_FROMHOST5_rst )
,.BRAM_FROMHOST5_addr( BRAM_FROMHOST5_addr )
,.BRAM_FROMHOST5_din( BRAM_FROMHOST5_din )
,.BRAM_FROMHOST5_dout( BRAM_FROMHOST5_dout )
,.BRAM_FROMHOST5_en( BRAM_FROMHOST5_en )
,.BRAM_FROMHOST5_we( BRAM_FROMHOST5_we )

,.BRAM_FROMHOST6_clk( BRAM_FROMHOST6_clk )
,.BRAM_FROMHOST6_rst( BRAM_FROMHOST6_rst )
,.BRAM_FROMHOST6_addr( BRAM_FROMHOST6_addr )
,.BRAM_FROMHOST6_din( BRAM_FROMHOST6_din )
,.BRAM_FROMHOST6_dout( BRAM_FROMHOST6_dout )
,.BRAM_FROMHOST6_en( BRAM_FROMHOST6_en )
,.BRAM_FROMHOST6_we( BRAM_FROMHOST6_we )

,.BRAM_FROMHOST7_clk( BRAM_FROMHOST7_clk )
,.BRAM_FROMHOST7_rst( BRAM_FROMHOST7_rst )
,.BRAM_FROMHOST7_addr( BRAM_FROMHOST7_addr )
,.BRAM_FROMHOST7_din( BRAM_FROMHOST7_din )
,.BRAM_FROMHOST7_dout( BRAM_FROMHOST7_dout )
,.BRAM_FROMHOST7_en( BRAM_FROMHOST7_en )
,.BRAM_FROMHOST7_we( BRAM_FROMHOST7_we )

,.BRAM_ACCBUF_clk( BRAM_ACCBUF_clk )
,.BRAM_ACCBUF_rst( BRAM_ACCBUF_rst )
,.BRAM_ACCBUF_addr( BRAM_ACCBUF_addr )
,.BRAM_ACCBUF_din( BRAM_ACCBUF_din )
,.BRAM_ACCBUF_dout( BRAM_ACCBUF_dout )
,.BRAM_ACCBUF_en( BRAM_ACCBUF_en )
,.BRAM_ACCBUF_we( BRAM_ACCBUF_we )

,.BRAM_COMMAND_clk( BRAM_COMMAND_clk )
,.BRAM_COMMAND_rst( BRAM_COMMAND_rst )
,.BRAM_COMMAND_addr( BRAM_COMMAND_addr )
,.BRAM_COMMAND_din( BRAM_COMMAND_din )
,.BRAM_COMMAND_dout( BRAM_COMMAND_dout )
,.BRAM_COMMAND_en( BRAM_COMMAND_en )
,.BRAM_COMMAND_we( BRAM_COMMAND_we )

,.clkadc2_300( clkadc2_300 )
,.clkadc2_600( clkadc2_600 )
,.DAC20_M_AXIS_ACLK( DAC20_M_AXIS_ACLK )
,.DAC20_M_AXIS_ARESETN( DAC20_M_AXIS_ARESETN )
,.DAC20_M_AXIS_TREADY( DAC20_M_AXIS_TREADY )
,.DAC20_M_AXIS_TVALID( DAC20_M_AXIS_TVALID )
,.DAC20_M_AXIS_TDATA( DAC20_M_AXIS_TDATA )
,.DAC20_M_AXIS_TSTRB( DAC20_M_AXIS_TSTRB )
,.DAC20_M_AXIS_TLAST( DAC20_M_AXIS_TLAST )
,.DAC22_M_AXIS_ACLK( DAC22_M_AXIS_ACLK )
,.DAC22_M_AXIS_ARESETN( DAC22_M_AXIS_ARESETN )
,.DAC22_M_AXIS_TREADY( DAC22_M_AXIS_TREADY )
,.DAC22_M_AXIS_TVALID( DAC22_M_AXIS_TVALID )
,.DAC22_M_AXIS_TDATA( DAC22_M_AXIS_TDATA )
,.DAC22_M_AXIS_TSTRB( DAC22_M_AXIS_TSTRB )
,.DAC22_M_AXIS_TLAST( DAC22_M_AXIS_TLAST )
,.clk_dac2( clk_dac2 )
,.DAC30_M_AXIS_ACLK( DAC30_M_AXIS_ACLK )
,.DAC30_M_AXIS_ARESETN( DAC30_M_AXIS_ARESETN )
,.DAC30_M_AXIS_TREADY( DAC30_M_AXIS_TREADY )
,.DAC30_M_AXIS_TVALID( DAC30_M_AXIS_TVALID )
,.DAC30_M_AXIS_TDATA( DAC30_M_AXIS_TDATA )
,.DAC30_M_AXIS_TSTRB( DAC30_M_AXIS_TSTRB )
,.DAC30_M_AXIS_TLAST( DAC30_M_AXIS_TLAST )
,.DAC32_M_AXIS_ACLK( DAC32_M_AXIS_ACLK )
,.DAC32_M_AXIS_ARESETN( DAC32_M_AXIS_ARESETN )
,.DAC32_M_AXIS_TREADY( DAC32_M_AXIS_TREADY )
,.DAC32_M_AXIS_TVALID( DAC32_M_AXIS_TVALID )
,.DAC32_M_AXIS_TDATA( DAC32_M_AXIS_TDATA )
,.DAC32_M_AXIS_TSTRB( DAC32_M_AXIS_TSTRB )
,.DAC32_M_AXIS_TLAST( DAC32_M_AXIS_TLAST )
,.clk_dac3( clk_dac3 )

,.ADC20_S_AXIS_ACLK( ADC20_S_AXIS_ACLK )
,.ADC20_S_AXIS_ARESETN( ADC20_S_AXIS_ARESETN )
,.ADC20_S_AXIS_TREADY( ADC20_S_AXIS_TREADY )
,.ADC20_S_AXIS_TVALID( ADC20_S_AXIS_TVALID )
,.ADC20_S_AXIS_TDATA( ADC20_S_AXIS_TDATA )
,.ADC20_S_AXIS_TSTRB( ADC20_S_AXIS_TSTRB )
,.ADC20_S_AXIS_TLAST( ADC20_S_AXIS_TLAST )
,.clk_adc2( clk_adc2 )
,.ADC21_S_AXIS_ACLK( ADC21_S_AXIS_ACLK )
,.ADC21_S_AXIS_ARESETN( ADC21_S_AXIS_ARESETN )
,.ADC21_S_AXIS_TREADY( ADC21_S_AXIS_TREADY )
,.ADC21_S_AXIS_TVALID( ADC21_S_AXIS_TVALID )
,.ADC21_S_AXIS_TDATA( ADC21_S_AXIS_TDATA )
,.ADC21_S_AXIS_TSTRB( ADC21_S_AXIS_TSTRB )
,.ADC21_S_AXIS_TLAST( ADC21_S_AXIS_TLAST )

,.cfgclk( cfgclk )
,.dspclk( dspclk )
