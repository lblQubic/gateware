ifbram acqbuf0_W
,ifbram acqbuf1_W
,ifbram command0_R
,ifbram command1_R
,ifbram command2_R
,ifbram command3_R
,ifbram command4_R
,ifbram command5_R
,ifbram command6_R
,ifbram command7_R
,ifbram qdrvfreq0_R
,ifbram qdrvfreq1_R
,ifbram qdrvfreq2_R
,ifbram qdrvfreq3_R
,ifbram qdrvfreq4_R
,ifbram qdrvfreq5_R
,ifbram qdrvfreq6_R
,ifbram qdrvfreq7_R
,ifbram rdrvfreq0_R
,ifbram rdrvfreq1_R
,ifbram rdrvfreq2_R
,ifbram rdrvfreq3_R
,ifbram rdrvfreq4_R
,ifbram rdrvfreq5_R
,ifbram rdrvfreq6_R
,ifbram rdrvfreq7_R
,ifbram dacmon0_W
,ifbram dacmon1_W
,ifbram dacmon2_W
,ifbram dacmon3_W
,ifbram qdrvenv0_R
,ifbram qdrvenv1_R
,ifbram qdrvenv2_R
,ifbram qdrvenv3_R
,ifbram qdrvenv4_R
,ifbram qdrvenv5_R
,ifbram qdrvenv6_R
,ifbram qdrvenv7_R
,ifbram rdloenv0_R
,ifbram rdloenv1_R
,ifbram rdloenv2_R
,ifbram rdloenv3_R
,ifbram rdloenv4_R
,ifbram rdloenv5_R
,ifbram rdloenv6_R
,ifbram rdloenv7_R
,ifbram rdrvenv0_R
,ifbram rdrvenv1_R
,ifbram rdrvenv2_R
,ifbram rdrvenv3_R
,ifbram rdrvenv4_R
,ifbram rdrvenv5_R
,ifbram rdrvenv6_R
,ifbram rdrvenv7_R
,ifbram accbuf0_W
,ifbram accbuf1_W
,ifbram accbuf2_W
,ifbram accbuf3_W
,ifbram accbuf4_W
,ifbram accbuf5_W
,ifbram accbuf6_W
,ifbram accbuf7_W
,ifbram rdlofreq0_R
,ifbram rdlofreq1_R
,ifbram rdlofreq2_R
,ifbram rdlofreq3_R
,ifbram rdlofreq4_R
,ifbram rdlofreq5_R
,ifbram rdlofreq6_R
,ifbram rdlofreq7_R
,ifbram sdbuf0_W
,ifbram sdbuf1_W
,ifbram sdbuf2_W
,ifbram sdbuf3_W
,ifbram sdbuf4_W
,ifbram sdbuf5_W
,ifbram sdbuf6_W
,ifbram sdbuf7_W