localparam INIT_acqbuf0="INIT_acqbuf0.mem";
localparam INIT_acqbuf1="INIT_acqbuf1.mem";
localparam INIT_command0="INIT_command0.mem";
localparam INIT_command1="INIT_command1.mem";
localparam INIT_command2="INIT_command2.mem";
localparam INIT_command3="INIT_command3.mem";
localparam INIT_command4="INIT_command4.mem";
localparam INIT_command5="INIT_command5.mem";
localparam INIT_command6="INIT_command6.mem";
localparam INIT_command7="INIT_command7.mem";
localparam INIT_qdrvfreq0="INIT_qdrvfreq0.mem";
localparam INIT_qdrvfreq1="INIT_qdrvfreq1.mem";
localparam INIT_qdrvfreq2="INIT_qdrvfreq2.mem";
localparam INIT_qdrvfreq3="INIT_qdrvfreq3.mem";
localparam INIT_qdrvfreq4="INIT_qdrvfreq4.mem";
localparam INIT_qdrvfreq5="INIT_qdrvfreq5.mem";
localparam INIT_qdrvfreq6="INIT_qdrvfreq6.mem";
localparam INIT_qdrvfreq7="INIT_qdrvfreq7.mem";
localparam INIT_rdrvfreq0="INIT_rdrvfreq0.mem";
localparam INIT_rdrvfreq1="INIT_rdrvfreq1.mem";
localparam INIT_rdrvfreq2="INIT_rdrvfreq2.mem";
localparam INIT_rdrvfreq3="INIT_rdrvfreq3.mem";
localparam INIT_rdrvfreq4="INIT_rdrvfreq4.mem";
localparam INIT_rdrvfreq5="INIT_rdrvfreq5.mem";
localparam INIT_rdrvfreq6="INIT_rdrvfreq6.mem";
localparam INIT_rdrvfreq7="INIT_rdrvfreq7.mem";
localparam INIT_dacmon0="INIT_dacmon0.mem";
localparam INIT_dacmon1="INIT_dacmon1.mem";
localparam INIT_dacmon2="INIT_dacmon2.mem";
localparam INIT_dacmon3="INIT_dacmon3.mem";
localparam INIT_qdrvenv0="INIT_qdrvenv0.mem";
localparam INIT_qdrvenv1="INIT_qdrvenv1.mem";
localparam INIT_qdrvenv2="INIT_qdrvenv2.mem";
localparam INIT_qdrvenv3="INIT_qdrvenv3.mem";
localparam INIT_qdrvenv4="INIT_qdrvenv4.mem";
localparam INIT_qdrvenv5="INIT_qdrvenv5.mem";
localparam INIT_qdrvenv6="INIT_qdrvenv6.mem";
localparam INIT_qdrvenv7="INIT_qdrvenv7.mem";
localparam INIT_rdloenv0="INIT_rdloenv0.mem";
localparam INIT_rdloenv1="INIT_rdloenv1.mem";
localparam INIT_rdloenv2="INIT_rdloenv2.mem";
localparam INIT_rdloenv3="INIT_rdloenv3.mem";
localparam INIT_rdloenv4="INIT_rdloenv4.mem";
localparam INIT_rdloenv5="INIT_rdloenv5.mem";
localparam INIT_rdloenv6="INIT_rdloenv6.mem";
localparam INIT_rdloenv7="INIT_rdloenv7.mem";
localparam INIT_rdrvenv0="INIT_rdrvenv0.mem";
localparam INIT_rdrvenv1="INIT_rdrvenv1.mem";
localparam INIT_rdrvenv2="INIT_rdrvenv2.mem";
localparam INIT_rdrvenv3="INIT_rdrvenv3.mem";
localparam INIT_rdrvenv4="INIT_rdrvenv4.mem";
localparam INIT_rdrvenv5="INIT_rdrvenv5.mem";
localparam INIT_rdrvenv6="INIT_rdrvenv6.mem";
localparam INIT_rdrvenv7="INIT_rdrvenv7.mem";
localparam INIT_accbuf0="INIT_accbuf0.mem";
localparam INIT_accbuf1="INIT_accbuf1.mem";
localparam INIT_accbuf2="INIT_accbuf2.mem";
localparam INIT_accbuf3="INIT_accbuf3.mem";
localparam INIT_accbuf4="INIT_accbuf4.mem";
localparam INIT_accbuf5="INIT_accbuf5.mem";
localparam INIT_accbuf6="INIT_accbuf6.mem";
localparam INIT_accbuf7="INIT_accbuf7.mem";
localparam INIT_rdlofreq0="INIT_rdlofreq0.mem";
localparam INIT_rdlofreq1="INIT_rdlofreq1.mem";
localparam INIT_rdlofreq2="INIT_rdlofreq2.mem";
localparam INIT_rdlofreq3="INIT_rdlofreq3.mem";
localparam INIT_rdlofreq4="INIT_rdlofreq4.mem";
localparam INIT_rdlofreq5="INIT_rdlofreq5.mem";
localparam INIT_rdlofreq6="INIT_rdlofreq6.mem";
localparam INIT_rdlofreq7="INIT_rdlofreq7.mem";
localparam INIT_sdbuf0="INIT_sdbuf0.mem";
localparam INIT_sdbuf1="INIT_sdbuf1.mem";
localparam INIT_sdbuf2="INIT_sdbuf2.mem";
localparam INIT_sdbuf3="INIT_sdbuf3.mem";
localparam INIT_sdbuf4="INIT_sdbuf4.mem";
localparam INIT_sdbuf5="INIT_sdbuf5.mem";
localparam INIT_sdbuf6="INIT_sdbuf6.mem";
localparam INIT_sdbuf7="INIT_sdbuf7.mem";