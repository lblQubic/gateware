module iladsp (input clk
,input [16-1:0] probe0
,input [16-1:0] probe1
,input [16-1:0] probe2
,input [16-1:0] probe3
,input [16-1:0] probe4
,input [16-1:0] probe5
,input [1-1:0] probe6
,input [4-1:0] probe7
,input [4-1:0] probe8
,input [1-1:0] probe9
,input [4-1:0] probe10
,input [4-1:0] probe11
,input [4-1:0] probe12
,input [4-1:0] probe13
,input [4-1:0] probe14
,input [4-1:0] probe15
,input [4-1:0] probe16
,input [4-1:0] probe17
,input [13-1:0] probe18
,input [64-1:0] probe19
,input [5-1:0] probe20
,input [5-1:0] probe21
,input [16-1:0] probe22
,input [16-1:0] probe23
,input [16-1:0] probe24
);
endmodule
