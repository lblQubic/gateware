.ACCBUF_R_ADDRWIDTH(ACCBUF_R_ADDRWIDTH),.ACCBUF_R_DATAWIDTH(ACCBUF_R_DATAWIDTH),.ACCBUF_W_ADDRWIDTH(ACCBUF_W_ADDRWIDTH),.ACCBUF_W_DATAWIDTH(ACCBUF_W_DATAWIDTH)
,.ACQBUF_R_ADDRWIDTH(ACQBUF_R_ADDRWIDTH),.ACQBUF_R_DATAWIDTH(ACQBUF_R_DATAWIDTH),.ACQBUF_W_ADDRWIDTH(ACQBUF_W_ADDRWIDTH),.ACQBUF_W_DATAWIDTH(ACQBUF_W_DATAWIDTH)
,.COMMAND_R_ADDRWIDTH(COMMAND_R_ADDRWIDTH),.COMMAND_R_DATAWIDTH(COMMAND_R_DATAWIDTH),.COMMAND_W_ADDRWIDTH(COMMAND_W_ADDRWIDTH),.COMMAND_W_DATAWIDTH(COMMAND_W_DATAWIDTH)
,.DACMON_R_ADDRWIDTH(DACMON_R_ADDRWIDTH),.DACMON_R_DATAWIDTH(DACMON_R_DATAWIDTH),.DACMON_W_ADDRWIDTH(DACMON_W_ADDRWIDTH),.DACMON_W_DATAWIDTH(DACMON_W_DATAWIDTH)
,.QDRVENV_R_ADDRWIDTH(QDRVENV_R_ADDRWIDTH),.QDRVENV_R_DATAWIDTH(QDRVENV_R_DATAWIDTH),.QDRVENV_W_ADDRWIDTH(QDRVENV_W_ADDRWIDTH),.QDRVENV_W_DATAWIDTH(QDRVENV_W_DATAWIDTH)
,.QDRVFREQ_R_ADDRWIDTH(QDRVFREQ_R_ADDRWIDTH),.QDRVFREQ_R_DATAWIDTH(QDRVFREQ_R_DATAWIDTH),.QDRVFREQ_W_ADDRWIDTH(QDRVFREQ_W_ADDRWIDTH),.QDRVFREQ_W_DATAWIDTH(QDRVFREQ_W_DATAWIDTH)
,.RDLOENV_R_ADDRWIDTH(RDLOENV_R_ADDRWIDTH),.RDLOENV_R_DATAWIDTH(RDLOENV_R_DATAWIDTH),.RDLOENV_W_ADDRWIDTH(RDLOENV_W_ADDRWIDTH),.RDLOENV_W_DATAWIDTH(RDLOENV_W_DATAWIDTH)
,.RDLOFREQ_R_ADDRWIDTH(RDLOFREQ_R_ADDRWIDTH),.RDLOFREQ_R_DATAWIDTH(RDLOFREQ_R_DATAWIDTH),.RDLOFREQ_W_ADDRWIDTH(RDLOFREQ_W_ADDRWIDTH),.RDLOFREQ_W_DATAWIDTH(RDLOFREQ_W_DATAWIDTH)
,.RDRVENV_R_ADDRWIDTH(RDRVENV_R_ADDRWIDTH),.RDRVENV_R_DATAWIDTH(RDRVENV_R_DATAWIDTH),.RDRVENV_W_ADDRWIDTH(RDRVENV_W_ADDRWIDTH),.RDRVENV_W_DATAWIDTH(RDRVENV_W_DATAWIDTH)
,.RDRVFREQ_R_ADDRWIDTH(RDRVFREQ_R_ADDRWIDTH),.RDRVFREQ_R_DATAWIDTH(RDRVFREQ_R_DATAWIDTH),.RDRVFREQ_W_ADDRWIDTH(RDRVFREQ_W_ADDRWIDTH),.RDRVFREQ_W_DATAWIDTH(RDRVFREQ_W_DATAWIDTH)